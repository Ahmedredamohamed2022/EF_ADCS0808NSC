magic
tech sky130A
magscale 1 2
timestamp 1686564671
<< checkpaint >>
rect -63314 -31298 45368 20457
<< nwell >>
rect -5990 13992 12994 14992
rect -5990 -25014 -4990 13992
rect 11994 9008 12994 13992
rect 11994 8008 39996 9008
rect 38996 -25014 39996 8008
rect -6002 -26014 39996 -25014
rect -5990 -26016 -4990 -26014
<< nsubdiff >>
rect -5914 14777 12894 14854
rect -5914 -25785 -5852 14777
rect -5274 14054 12168 14199
rect -5274 -25098 -5114 14054
rect 12094 8351 12168 14054
rect 12746 8948 12894 14777
rect 12746 8861 39904 8948
rect 12094 8148 39232 8351
rect 39104 -25098 39232 8148
rect -5274 -25207 39232 -25098
rect 39810 -25785 39904 8861
rect -5914 -25856 39904 -25785
rect -5904 -25898 39904 -25856
<< nsubdiffcont >>
rect -5852 14199 12746 14777
rect -5852 -25207 -5274 14199
rect 12168 8861 12746 14199
rect 12168 8351 39810 8861
rect 39232 -25207 39810 8351
rect -5852 -25785 39810 -25207
<< locali >>
rect -5926 14781 12906 14854
rect -5926 14777 -5823 14781
rect 12715 14777 12906 14781
rect -5926 -25785 -5852 14777
rect -5274 14054 12168 14199
rect -5274 -25056 -5126 14054
rect 12106 8351 12168 14054
rect 12746 8938 12906 14777
rect 12746 8877 39904 8938
rect 39787 8861 39904 8877
rect 12106 8339 12177 8351
rect 12106 8138 39232 8339
rect 39104 -25056 39232 8138
rect -5274 -25207 39232 -25056
rect 39810 -25785 39904 8861
rect -5926 -25789 -5823 -25785
rect 39787 -25789 39904 -25785
rect -5926 -25856 39904 -25789
<< viali >>
rect -5823 14777 12715 14781
rect -5823 14243 12715 14777
rect -5823 -25251 -5285 14243
rect 12177 8877 12715 14243
rect 12177 8861 12746 8877
rect 12746 8861 39787 8877
rect 12177 8351 39787 8861
rect 12177 8339 39232 8351
rect 39232 8339 39787 8351
rect 39249 -25251 39787 8339
rect -5823 -25785 39787 -25251
rect -5823 -25789 39787 -25785
<< metal1 >>
rect -6000 14781 12990 14968
rect -6000 -25789 -5823 14781
rect -5285 13968 12177 14243
rect -5285 -25016 -5000 13968
rect 11990 8339 12177 13968
rect 12715 9016 12990 14781
rect 12715 8877 39996 9016
rect 11990 8016 39249 8339
rect 23008 4923 23600 5002
rect 23008 4487 23061 4923
rect 23497 4487 23600 4923
rect 23008 4404 23600 4487
rect 24664 4971 25250 5042
rect 24664 4535 24717 4971
rect 25153 4535 25250 4971
rect 24664 4456 25250 4535
rect 26416 4973 27002 5044
rect 26416 4537 26469 4973
rect 26905 4537 27002 4973
rect 26416 4458 27002 4537
rect 28066 4971 28652 5042
rect 28066 4535 28119 4971
rect 28555 4535 28652 4971
rect 28066 4456 28652 4535
rect 29590 4959 30176 5030
rect 29590 4523 29643 4959
rect 30079 4523 30176 4959
rect 29590 4444 30176 4523
rect 31280 4999 31866 5070
rect 31280 4563 31333 4999
rect 31769 4563 31866 4999
rect 31280 4484 31866 4563
rect 32866 4999 33452 5070
rect 32866 4563 32919 4999
rect 33355 4563 33452 4999
rect 32866 4484 33452 4563
rect 34466 4969 35052 5040
rect 34466 4533 34519 4969
rect 34955 4533 35052 4969
rect 34466 4454 35052 4533
rect 16974 1906 17974 1978
rect 16974 1214 17051 1906
rect 17807 1746 17974 1906
rect 17807 1384 21924 1746
rect 17807 1214 17974 1384
rect 16974 1038 17974 1214
rect 4396 -2180 4802 -1998
rect 4396 -2360 4470 -2180
rect 4714 -2360 4802 -2180
rect 4396 -2400 4802 -2360
rect 4396 -2518 4804 -2400
rect 4396 -2520 4802 -2518
rect 10764 -10594 11086 -10540
rect 10764 -10966 10794 -10594
rect 11038 -10966 11086 -10594
rect 10764 -11006 11086 -10966
rect 94 -21686 490 -21646
rect -688 -21804 -342 -21794
rect -688 -22036 -200 -21804
rect -688 -22664 -599 -22036
rect -291 -22664 -200 -22036
rect 94 -22122 162 -21686
rect 406 -22122 490 -21686
rect 2000 -21683 3122 -21604
rect 2000 -21927 2090 -21683
rect 3038 -21927 3122 -21683
rect 4076 -21672 4296 -21608
rect 2000 -22006 3122 -21927
rect 3254 -21871 3992 -21728
rect 94 -22200 490 -22122
rect 3254 -22499 3349 -21871
rect 3913 -22499 3992 -21871
rect 4076 -22300 4099 -21672
rect 4279 -22300 4296 -21672
rect 4076 -22364 4296 -22300
rect 4430 -21762 4628 -21694
rect 4430 -22326 4471 -21762
rect 4587 -22326 4628 -21762
rect 4430 -22392 4628 -22326
rect 3254 -22508 3992 -22499
rect -688 -22776 -200 -22664
rect -682 -22782 -200 -22776
rect 38996 -25016 39249 8016
rect -5285 -25251 39249 -25016
rect 39787 -25789 39996 8877
rect -6000 -25994 39996 -25789
rect -5990 -26016 39996 -25994
<< via1 >>
rect 23061 4487 23497 4923
rect 24717 4535 25153 4971
rect 26469 4537 26905 4973
rect 28119 4535 28555 4971
rect 29643 4523 30079 4959
rect 31333 4563 31769 4999
rect 32919 4563 33355 4999
rect 34519 4533 34955 4969
rect 17051 1214 17807 1906
rect 4470 -2360 4714 -2180
rect 10794 -10966 11038 -10594
rect -599 -22664 -291 -22036
rect 162 -22122 406 -21686
rect 2090 -21927 3038 -21683
rect 3349 -22499 3913 -21871
rect 4099 -22300 4279 -21672
rect 4471 -22326 4587 -21762
<< metal2 >>
rect -4004 12478 11020 13502
rect -4004 2865 -2980 12478
rect 8044 11625 9026 11834
rect 8044 11300 8152 11625
rect 4190 11200 4794 11244
rect 4190 11064 4254 11200
rect 4710 11064 4794 11200
rect 1974 10963 3614 11054
rect 4190 10996 4794 11064
rect 1974 10507 2234 10963
rect 3490 10507 3614 10963
rect 1974 10352 3614 10507
rect 4282 10200 4366 10996
rect 8030 9569 8152 11300
rect 8848 10994 9026 11625
rect 8848 9569 8998 10994
rect 8030 8940 8998 9569
rect 9996 6974 11020 12478
rect 9996 5950 38012 6974
rect 20392 5682 20784 5760
rect 20366 5582 20784 5682
rect 20366 3766 20479 5582
rect 20695 3766 20784 5582
rect 20916 5514 21226 5642
rect 20916 3858 20978 5514
rect 21194 3858 21226 5514
rect 23008 4923 23600 5002
rect 23008 4893 23061 4923
rect 23497 4893 23600 4923
rect 23008 4517 23051 4893
rect 23507 4517 23600 4893
rect 23008 4487 23061 4517
rect 23497 4487 23600 4517
rect 23008 4404 23600 4487
rect 24664 4971 25250 5042
rect 24664 4941 24717 4971
rect 25153 4941 25250 4971
rect 24664 4565 24707 4941
rect 25163 4565 25250 4941
rect 24664 4535 24717 4565
rect 25153 4535 25250 4565
rect 24664 4456 25250 4535
rect 26416 4973 27002 5044
rect 26416 4943 26469 4973
rect 26905 4943 27002 4973
rect 26416 4567 26459 4943
rect 26915 4567 27002 4943
rect 26416 4537 26469 4567
rect 26905 4537 27002 4567
rect 26416 4458 27002 4537
rect 28066 4971 28652 5042
rect 28066 4941 28119 4971
rect 28555 4941 28652 4971
rect 28066 4565 28109 4941
rect 28565 4565 28652 4941
rect 28066 4535 28119 4565
rect 28555 4535 28652 4565
rect 28066 4456 28652 4535
rect 29590 4959 30176 5030
rect 29590 4929 29643 4959
rect 30079 4929 30176 4959
rect 29590 4553 29633 4929
rect 30089 4553 30176 4929
rect 29590 4523 29643 4553
rect 30079 4523 30176 4553
rect 29590 4444 30176 4523
rect 31280 4999 31866 5070
rect 31280 4969 31333 4999
rect 31769 4969 31866 4999
rect 31280 4593 31323 4969
rect 31779 4593 31866 4969
rect 31280 4563 31333 4593
rect 31769 4563 31866 4593
rect 31280 4484 31866 4563
rect 32866 4999 33452 5070
rect 32866 4969 32919 4999
rect 33355 4969 33452 4999
rect 32866 4593 32909 4969
rect 33365 4593 33452 4969
rect 32866 4563 32919 4593
rect 33355 4563 33452 4593
rect 32866 4484 33452 4563
rect 34466 4969 35052 5040
rect 34466 4939 34519 4969
rect 34955 4939 35052 4969
rect 34466 4563 34509 4939
rect 34965 4563 35052 4939
rect 34466 4533 34519 4563
rect 34955 4533 35052 4563
rect 34466 4454 35052 4533
rect 20916 3768 21226 3858
rect 20366 3606 20784 3766
rect 20366 3584 20770 3606
rect -4004 1929 -3938 2865
rect -3082 1929 -2980 2865
rect -4004 -22986 -2980 1929
rect 16974 1908 17974 1978
rect 16974 1906 17081 1908
rect 17777 1906 17974 1908
rect 16974 1214 17051 1906
rect 17807 1214 17974 1906
rect 16974 1212 17081 1214
rect 17777 1212 17974 1214
rect 16974 1038 17974 1212
rect 5364 -1814 5448 -1002
rect 5594 -1734 5694 -832
rect 4386 -1877 5472 -1814
rect 4386 -2093 5034 -1877
rect 5410 -2093 5472 -1877
rect 4386 -2154 5472 -2093
rect 5594 -1899 7066 -1734
rect 4396 -2157 4802 -2154
rect 4396 -2373 4444 -2157
rect 4740 -2373 4802 -2157
rect 5594 -2195 6137 -1899
rect 6833 -2195 7066 -1899
rect 5594 -2286 7066 -2195
rect 5596 -2316 7066 -2286
rect 4396 -2400 4802 -2373
rect 4396 -2518 4804 -2400
rect 4396 -2520 4802 -2518
rect 10764 -10592 11086 -10540
rect 10764 -10594 10808 -10592
rect 11024 -10594 11086 -10592
rect 10764 -10966 10794 -10594
rect 11038 -10966 11086 -10594
rect 10764 -10968 10808 -10966
rect 11024 -10968 11086 -10966
rect 10764 -11006 11086 -10968
rect 36988 -20618 38012 5950
rect 36988 -20834 37080 -20618
rect 37936 -20834 38012 -20618
rect 94 -21686 490 -21646
rect -682 -22036 -200 -21804
rect -682 -22664 -599 -22036
rect -291 -22664 -200 -22036
rect 94 -22122 162 -21686
rect 406 -22122 490 -21686
rect 2000 -21683 3122 -21604
rect 2000 -21927 2090 -21683
rect 3038 -21927 3122 -21683
rect 4076 -21672 4296 -21608
rect 2000 -22006 3122 -21927
rect 3254 -21871 3992 -21728
rect 94 -22200 490 -22122
rect 3254 -22499 3349 -21871
rect 3913 -22499 3992 -21871
rect 4076 -22300 4099 -21672
rect 4279 -22300 4296 -21672
rect 4076 -22364 4296 -22300
rect 4430 -21762 4628 -21694
rect 4430 -21776 4471 -21762
rect 4587 -21776 4628 -21762
rect 4430 -22312 4461 -21776
rect 4597 -22312 4628 -21776
rect 4430 -22326 4471 -22312
rect 4587 -22326 4628 -22312
rect 4430 -22392 4628 -22326
rect 3254 -22508 3992 -22499
rect -682 -22782 -200 -22664
rect 36988 -22986 38012 -20834
rect -4040 -23078 38012 -22986
rect -4040 -23854 -1888 -23078
rect -1032 -23854 38012 -23078
rect -4040 -24010 38012 -23854
<< via2 >>
rect 4254 11064 4710 11200
rect 2234 10507 3490 10963
rect 8152 9569 8848 11625
rect 20479 3766 20695 5582
rect 20978 3858 21194 5514
rect 23051 4517 23061 4893
rect 23061 4517 23497 4893
rect 23497 4517 23507 4893
rect 24707 4565 24717 4941
rect 24717 4565 25153 4941
rect 25153 4565 25163 4941
rect 26459 4567 26469 4943
rect 26469 4567 26905 4943
rect 26905 4567 26915 4943
rect 28109 4565 28119 4941
rect 28119 4565 28555 4941
rect 28555 4565 28565 4941
rect 29633 4553 29643 4929
rect 29643 4553 30079 4929
rect 30079 4553 30089 4929
rect 31323 4593 31333 4969
rect 31333 4593 31769 4969
rect 31769 4593 31779 4969
rect 32909 4593 32919 4969
rect 32919 4593 33355 4969
rect 33355 4593 33365 4969
rect 34509 4563 34519 4939
rect 34519 4563 34955 4939
rect 34955 4563 34965 4939
rect -3938 1929 -3082 2865
rect 17081 1906 17777 1908
rect 17081 1214 17777 1906
rect 17081 1212 17777 1214
rect 5034 -2093 5410 -1877
rect 4444 -2180 4740 -2157
rect 4444 -2360 4470 -2180
rect 4470 -2360 4714 -2180
rect 4714 -2360 4740 -2180
rect 4444 -2373 4740 -2360
rect 6137 -2195 6833 -1899
rect 10808 -10594 11024 -10592
rect 10808 -10966 11024 -10594
rect 10808 -10968 11024 -10966
rect 37080 -20834 37936 -20618
rect -593 -22658 -297 -22042
rect 176 -22092 392 -21716
rect 2096 -21913 3032 -21697
rect 3363 -22493 3899 -21877
rect 4121 -22294 4257 -21678
rect 4461 -22312 4471 -21776
rect 4471 -22312 4587 -21776
rect 4587 -22312 4597 -21776
rect -1888 -23854 -1032 -23078
<< metal3 >>
rect -61812 18885 -60702 19102
rect -61812 18181 -61713 18885
rect -60849 18181 -60702 18885
rect -61812 -29165 -60702 18181
rect -61812 -29869 -61789 -29165
rect -60925 -29869 -60702 -29165
rect -61812 -29970 -60702 -29869
rect -60112 16889 -59002 19102
rect -60112 16185 -59959 16889
rect -59095 16185 -59002 16889
rect -60112 -27151 -59002 16185
rect -9890 18865 -8952 19056
rect -9890 18161 -9754 18865
rect -9130 18161 -8952 18865
rect -9890 15440 -8952 18161
rect -8098 17084 -7012 17180
rect -8098 16060 -7771 17084
rect -7147 16060 -7012 17084
rect -8098 15440 -7012 16060
rect -9898 11003 -8870 15440
rect -8098 14472 -6972 15440
rect -9898 10379 -9730 11003
rect -9026 10379 -8870 11003
rect -9898 6138 -8870 10379
rect -9898 2794 -9737 6138
rect -9033 2794 -8870 6138
rect -9898 -10702 -8870 2794
rect -9898 -11406 -9777 -10702
rect -8993 -11406 -8870 -10702
rect -57264 -12178 -56186 -12064
rect -57246 -12550 -56168 -12436
rect -57214 -12928 -56136 -12814
rect -57216 -13308 -56138 -13194
rect -57342 -16646 -56264 -16532
rect -57344 -19358 -56266 -19244
rect -57324 -21934 -56246 -21820
rect -57374 -25348 -56296 -25234
rect -57372 -25738 -56294 -25624
rect -57352 -26098 -56274 -25984
rect -57344 -26484 -56266 -26370
rect -60112 -27855 -60015 -27151
rect -59151 -27855 -59002 -27151
rect -60112 -29970 -59002 -27855
rect -9898 -29134 -8870 -11406
rect -8000 12085 -6972 14472
rect -8000 11541 -7936 12085
rect -7072 11541 -6972 12085
rect -8000 -27120 -6972 11541
rect -5992 14968 -5002 14998
rect -5992 14104 -5787 14968
rect -5163 14104 -5002 14968
rect -5992 560 -5002 14104
rect 20922 12949 21262 13092
rect 20922 12085 20976 12949
rect 21200 12085 21262 12949
rect 8044 11629 9026 11834
rect 8044 11625 8188 11629
rect 8812 11625 9026 11629
rect 8044 11300 8152 11625
rect 4190 11204 4794 11244
rect 4190 11200 4290 11204
rect 4674 11200 4794 11204
rect 4190 11064 4254 11200
rect 4710 11064 4794 11200
rect 4190 11060 4290 11064
rect 4674 11060 4794 11064
rect 1974 10967 3614 11054
rect 4190 10996 4794 11060
rect 1974 10503 2230 10967
rect 3494 10503 3614 10967
rect 1974 10352 3614 10503
rect 8030 9569 8152 11300
rect 8848 10994 9026 11625
rect 8848 9569 8998 10994
rect 8030 9565 8188 9569
rect 8812 9565 8998 9569
rect 8030 8940 8998 9565
rect 20394 10956 20784 11060
rect 20394 10012 20417 10956
rect 20721 10012 20784 10956
rect 20394 5682 20784 10012
rect 20366 5582 20784 5682
rect 20922 5642 21262 12085
rect 42914 12878 43938 13042
rect 42914 12014 43085 12878
rect 43789 12014 43938 12878
rect 40910 10956 41976 11016
rect 40910 10012 41154 10956
rect 41858 10012 41976 10956
rect 20366 3766 20479 5582
rect 20695 3766 20784 5582
rect 20916 5514 21262 5642
rect 20916 3858 20978 5514
rect 21194 3858 21262 5514
rect 38884 9018 39992 9098
rect 38884 8154 39192 9018
rect 39896 8154 39992 9018
rect 23008 4897 23600 5002
rect 23008 4513 23047 4897
rect 23511 4513 23600 4897
rect 23008 4404 23600 4513
rect 24664 4945 25250 5042
rect 24664 4561 24703 4945
rect 25167 4561 25250 4945
rect 24664 4456 25250 4561
rect 26416 4947 27002 5044
rect 26416 4563 26455 4947
rect 26919 4563 27002 4947
rect 26416 4458 27002 4563
rect 28066 4945 28652 5042
rect 28066 4561 28105 4945
rect 28569 4561 28652 4945
rect 28066 4456 28652 4561
rect 29590 4933 30176 5030
rect 29590 4549 29629 4933
rect 30093 4549 30176 4933
rect 29590 4444 30176 4549
rect 31280 4973 31866 5070
rect 31280 4589 31319 4973
rect 31783 4589 31866 4973
rect 31280 4484 31866 4589
rect 32866 4973 33452 5070
rect 32866 4589 32905 4973
rect 33369 4589 33452 4973
rect 32866 4484 33452 4589
rect 34466 4943 35052 5040
rect 34466 4559 34505 4943
rect 34969 4559 35052 4943
rect 34466 4454 35052 4559
rect 20916 3768 21262 3858
rect 20366 3628 20784 3766
rect 20922 3744 21262 3768
rect 20366 3584 20770 3628
rect -3990 2869 -3002 2938
rect -3990 2865 -3902 2869
rect -3118 2865 -3002 2869
rect -3990 1929 -3938 2865
rect -3082 1929 -3002 2865
rect 9634 2134 10198 2142
rect -3990 1925 -3902 1929
rect -3118 1925 -3002 1929
rect -3990 1848 -3002 1925
rect 9468 1925 10218 2134
rect 9468 1061 9599 1925
rect 10143 1061 10218 1925
rect 9468 956 10218 1061
rect 16974 1912 17974 1978
rect 16974 1208 17077 1912
rect 17781 1208 17974 1912
rect 16974 1038 17974 1208
rect -5992 -384 -5825 560
rect -5121 -384 -5002 560
rect -5992 -25122 -5002 -384
rect 4386 -1873 5472 -1814
rect 4386 -2075 5030 -1873
rect 4386 -2154 4440 -2075
rect 4396 -2379 4440 -2154
rect 4744 -2097 5030 -2075
rect 5414 -2097 5472 -1873
rect 4744 -2154 5472 -2097
rect 5596 -1895 7066 -1734
rect 4744 -2379 4802 -2154
rect 5596 -2199 6133 -1895
rect 6837 -2199 7066 -1895
rect 5596 -2316 7066 -2199
rect 4396 -2514 4802 -2379
rect 94 -21712 490 -21646
rect -682 -22038 -200 -21804
rect -682 -22570 -597 -22038
rect -700 -22662 -597 -22570
rect -293 -22662 -200 -22038
rect 94 -22096 172 -21712
rect 396 -22096 490 -21712
rect 2000 -21693 3122 -21604
rect 2000 -21917 2092 -21693
rect 3036 -21917 3122 -21693
rect 4076 -21674 4296 -21608
rect 2000 -22006 3122 -21917
rect 3254 -21873 3992 -21728
rect 94 -22200 490 -22096
rect -700 -22782 -200 -22662
rect -1994 -23074 -926 -22958
rect -1994 -23858 -1892 -23074
rect -1028 -23858 -926 -23074
rect -1994 -23996 -926 -23858
rect -5992 -25906 -5863 -25122
rect -5079 -25906 -5002 -25122
rect -5992 -25986 -5002 -25906
rect -8000 -27904 -7903 -27120
rect -7119 -27904 -6972 -27120
rect -8000 -28014 -6972 -27904
rect -700 -28982 -214 -22782
rect 2026 -26982 3096 -22006
rect 3254 -22497 3359 -21873
rect 3903 -22497 3992 -21873
rect 4076 -22298 4117 -21674
rect 4261 -22298 4296 -21674
rect 4076 -22364 4296 -22298
rect 4430 -21772 4628 -21694
rect 4430 -22316 4457 -21772
rect 4601 -22316 4628 -21772
rect 4430 -22392 4628 -22316
rect 9634 -21987 10198 956
rect 10776 -1802 11046 -1696
rect 10776 -2266 10810 -1802
rect 11034 -2266 11046 -1802
rect 10776 -10540 11046 -2266
rect 35560 -2109 36264 -2042
rect 35560 -2413 35598 -2109
rect 36222 -2413 36264 -2109
rect 35560 -2508 36264 -2413
rect 38884 -2117 39992 8154
rect 38884 -2421 39125 -2117
rect 39909 -2421 39992 -2117
rect 35576 -2647 36518 -2600
rect 35576 -2791 35697 -2647
rect 36401 -2791 36518 -2647
rect 35576 -2832 36518 -2791
rect 10764 -10592 11086 -10540
rect 10764 -10968 10808 -10592
rect 11024 -10968 11086 -10592
rect 10764 -11006 11086 -10968
rect 35580 -20279 36510 -20240
rect 35580 -20423 35676 -20279
rect 36460 -20423 36510 -20279
rect 35580 -20466 36510 -20423
rect 35624 -20618 38002 -20532
rect 35624 -20834 37080 -20618
rect 37936 -20834 38002 -20618
rect 35624 -20900 38002 -20834
rect 9634 -22291 9670 -21987
rect 10134 -22291 10198 -21987
rect 9634 -22412 10198 -22291
rect 3254 -22508 3992 -22497
rect 3270 -22796 3980 -22508
rect 3270 -24332 3963 -22796
rect 3270 -25025 3980 -24332
rect 3270 -25889 3381 -25025
rect 3925 -25889 3980 -25025
rect 38884 -24969 39992 -2421
rect 38884 -25593 39169 -24969
rect 39793 -25593 39992 -24969
rect 38884 -25836 39992 -25593
rect 3270 -25978 3980 -25889
rect 1986 -27117 3096 -26982
rect 1986 -27901 2131 -27117
rect 2915 -27810 3096 -27117
rect 40910 -27054 41976 10012
rect 2915 -27901 3074 -27810
rect 1986 -28044 3074 -27901
rect 40910 -27838 41059 -27054
rect 41763 -27838 41976 -27054
rect 40910 -27990 41976 -27838
rect -9898 -29918 -9761 -29134
rect -8977 -29918 -8870 -29134
rect -9898 -30030 -8870 -29918
rect -1036 -29124 68 -28982
rect -1036 -29828 -810 -29124
rect -186 -29828 68 -29124
rect -1036 -30038 68 -29828
rect 42914 -29151 43938 12014
rect 42914 -29855 43199 -29151
rect 43823 -29855 43938 -29151
rect 42914 -30016 43938 -29855
<< via3 >>
rect -61713 18181 -60849 18885
rect -61789 -29869 -60925 -29165
rect -59959 16185 -59095 16889
rect -9754 18161 -9130 18865
rect -7771 16060 -7147 17084
rect -9730 10379 -9026 11003
rect -9737 2794 -9033 6138
rect -9777 -11406 -8993 -10702
rect -60015 -27855 -59151 -27151
rect -7936 11541 -7072 12085
rect -5787 14104 -5163 14968
rect 20976 12085 21200 12949
rect 8188 11625 8812 11629
rect 4290 11200 4674 11204
rect 4290 11064 4674 11200
rect 4290 11060 4674 11064
rect 2230 10963 3494 10967
rect 2230 10507 2234 10963
rect 2234 10507 3490 10963
rect 3490 10507 3494 10963
rect 2230 10503 3494 10507
rect 8188 9569 8812 11625
rect 8188 9565 8812 9569
rect 20417 10012 20721 10956
rect 43085 12014 43789 12878
rect 41154 10012 41858 10956
rect 39192 8154 39896 9018
rect 23047 4893 23511 4897
rect 23047 4517 23051 4893
rect 23051 4517 23507 4893
rect 23507 4517 23511 4893
rect 23047 4513 23511 4517
rect 24703 4941 25167 4945
rect 24703 4565 24707 4941
rect 24707 4565 25163 4941
rect 25163 4565 25167 4941
rect 24703 4561 25167 4565
rect 26455 4943 26919 4947
rect 26455 4567 26459 4943
rect 26459 4567 26915 4943
rect 26915 4567 26919 4943
rect 26455 4563 26919 4567
rect 28105 4941 28569 4945
rect 28105 4565 28109 4941
rect 28109 4565 28565 4941
rect 28565 4565 28569 4941
rect 28105 4561 28569 4565
rect 29629 4929 30093 4933
rect 29629 4553 29633 4929
rect 29633 4553 30089 4929
rect 30089 4553 30093 4929
rect 29629 4549 30093 4553
rect 31319 4969 31783 4973
rect 31319 4593 31323 4969
rect 31323 4593 31779 4969
rect 31779 4593 31783 4969
rect 31319 4589 31783 4593
rect 32905 4969 33369 4973
rect 32905 4593 32909 4969
rect 32909 4593 33365 4969
rect 33365 4593 33369 4969
rect 32905 4589 33369 4593
rect 34505 4939 34969 4943
rect 34505 4563 34509 4939
rect 34509 4563 34965 4939
rect 34965 4563 34969 4939
rect 34505 4559 34969 4563
rect -3902 2865 -3118 2869
rect -3902 1929 -3118 2865
rect -3902 1925 -3118 1929
rect 9599 1061 10143 1925
rect 17077 1908 17781 1912
rect 17077 1212 17081 1908
rect 17081 1212 17777 1908
rect 17777 1212 17781 1908
rect 17077 1208 17781 1212
rect -5825 -384 -5121 560
rect 5030 -1877 5414 -1873
rect 4440 -2157 4744 -2075
rect 5030 -2093 5034 -1877
rect 5034 -2093 5410 -1877
rect 5410 -2093 5414 -1877
rect 5030 -2097 5414 -2093
rect 4440 -2373 4444 -2157
rect 4444 -2373 4740 -2157
rect 4740 -2373 4744 -2157
rect 4440 -2379 4744 -2373
rect 6133 -1899 6837 -1895
rect 6133 -2195 6137 -1899
rect 6137 -2195 6833 -1899
rect 6833 -2195 6837 -1899
rect 6133 -2199 6837 -2195
rect -597 -22042 -293 -22038
rect -597 -22658 -593 -22042
rect -593 -22658 -297 -22042
rect -297 -22658 -293 -22042
rect -597 -22662 -293 -22658
rect 172 -21716 396 -21712
rect 172 -22092 176 -21716
rect 176 -22092 392 -21716
rect 392 -22092 396 -21716
rect 172 -22096 396 -22092
rect 2092 -21697 3036 -21693
rect 2092 -21913 2096 -21697
rect 2096 -21913 3032 -21697
rect 3032 -21913 3036 -21697
rect 2092 -21917 3036 -21913
rect -1892 -23078 -1028 -23074
rect -1892 -23854 -1888 -23078
rect -1888 -23854 -1032 -23078
rect -1032 -23854 -1028 -23078
rect -1892 -23858 -1028 -23854
rect -5863 -25906 -5079 -25122
rect -7903 -27904 -7119 -27120
rect 3359 -21877 3903 -21873
rect 3359 -22493 3363 -21877
rect 3363 -22493 3899 -21877
rect 3899 -22493 3903 -21877
rect 3359 -22497 3903 -22493
rect 4117 -21678 4261 -21674
rect 4117 -22294 4121 -21678
rect 4121 -22294 4257 -21678
rect 4257 -22294 4261 -21678
rect 4117 -22298 4261 -22294
rect 4457 -21776 4601 -21772
rect 4457 -22312 4461 -21776
rect 4461 -22312 4597 -21776
rect 4597 -22312 4601 -21776
rect 4457 -22316 4601 -22312
rect 10810 -2266 11034 -1802
rect 35598 -2413 36222 -2109
rect 39125 -2421 39909 -2117
rect 35697 -2791 36401 -2647
rect 35676 -20423 36460 -20279
rect 9670 -22291 10134 -21987
rect 3381 -25889 3925 -25025
rect 39169 -25593 39793 -24969
rect 2131 -27901 2915 -27117
rect 41059 -27838 41763 -27054
rect -9761 -29918 -8977 -29134
rect -810 -29828 -186 -29124
rect 43199 -29855 43823 -29151
<< metal4 >>
rect 15936 19014 16982 19078
rect -62054 18885 16982 19014
rect -62054 18181 -61713 18885
rect -60849 18865 16982 18885
rect -60849 18181 -9754 18865
rect -62054 18161 -9754 18181
rect -9130 18161 16982 18865
rect -62054 18034 16982 18161
rect -62054 17084 14934 17202
rect -62054 16889 -7771 17084
rect -62054 16185 -59959 16889
rect -59095 16185 -7771 16889
rect -62054 16060 -7771 16185
rect -7147 17052 14934 17084
rect -7147 16060 14976 17052
rect -62054 15964 14976 16060
rect -5966 15068 13056 15090
rect -5966 14968 13120 15068
rect -5966 14104 -5787 14968
rect -5163 14104 13120 14968
rect -5966 13982 13120 14104
rect -3244 12190 9002 12202
rect -8094 12085 9002 12190
rect -8094 11541 -7936 12085
rect -7072 11924 9002 12085
rect -7072 11629 9026 11924
rect -7072 11541 8188 11629
rect -8094 11450 8188 11541
rect -7924 11436 8188 11450
rect 8044 11300 8188 11436
rect 4190 11204 4794 11244
rect -10044 11054 2670 11088
rect 4190 11060 4290 11204
rect 4674 11060 4794 11204
rect -10044 11003 3614 11054
rect -10044 10379 -9730 11003
rect -9026 10967 3614 11003
rect 4190 10996 4794 11060
rect -9026 10503 2230 10967
rect 3494 10503 3614 10967
rect -9026 10379 3614 10503
rect -10044 10352 3614 10379
rect -10044 10336 2670 10352
rect 8030 9565 8188 11300
rect 8812 10994 9026 11629
rect 8812 9565 8998 10994
rect 8030 8940 8998 9565
rect 11948 9140 13120 13982
rect 13974 11102 14976 15964
rect 15936 13106 16982 18034
rect 15936 12949 44108 13106
rect 15936 12085 20976 12949
rect 21200 12878 44108 12949
rect 21200 12085 43085 12878
rect 15936 12040 43085 12085
rect 15978 12014 43085 12040
rect 43789 12014 44108 12878
rect 15978 11976 44108 12014
rect 13952 10956 41954 11102
rect 13952 10012 20417 10956
rect 20721 10012 41154 10956
rect 41858 10012 41954 10956
rect 13952 9908 41954 10012
rect 11948 9018 40034 9140
rect 11948 8202 39192 9018
rect 12012 8154 39192 8202
rect 39896 8154 40034 9018
rect 12012 8074 40034 8154
rect -9940 6138 -8912 6302
rect -9940 4649 -9737 6138
rect -21792 3689 -9737 4649
rect -9940 2794 -9737 3689
rect -9033 4649 -8912 6138
rect 23008 4897 23600 5002
rect -9033 3689 -8892 4649
rect 23008 4513 23047 4897
rect 23511 4513 23600 4897
rect 23008 4404 23600 4513
rect 24664 4945 25250 5042
rect 24664 4561 24703 4945
rect 25167 4561 25250 4945
rect 24664 4456 25250 4561
rect 26416 4947 27002 5044
rect 26416 4563 26455 4947
rect 26919 4563 27002 4947
rect 26416 4458 27002 4563
rect 28066 4945 28652 5042
rect 28066 4561 28105 4945
rect 28569 4561 28652 4945
rect 28066 4456 28652 4561
rect 29590 4933 30176 5030
rect 29590 4549 29629 4933
rect 30093 4549 30176 4933
rect 29590 4444 30176 4549
rect 31280 4973 31866 5070
rect 31280 4589 31319 4973
rect 31783 4589 31866 4973
rect 31280 4484 31866 4589
rect 32866 4973 33452 5070
rect 32866 4589 32905 4973
rect 33369 4589 33452 4973
rect 32866 4484 33452 4589
rect 34466 4943 35052 5040
rect 34466 4559 34505 4943
rect 34969 4559 35052 4943
rect 34466 4454 35052 4559
rect -9033 2794 -8912 3689
rect -9940 2412 -8912 2794
rect -3998 2869 -830 2944
rect -3998 1925 -3902 2869
rect -3118 1925 -830 2869
rect -3998 1816 -830 1925
rect 9468 1994 10218 2134
rect 9468 1978 17958 1994
rect 9468 1925 17974 1978
rect 9468 1061 9599 1925
rect 10143 1912 17974 1925
rect 10143 1208 17077 1912
rect 17781 1208 17974 1912
rect 10143 1061 17974 1208
rect 9468 1038 17974 1061
rect 9468 956 17958 1038
rect 9536 948 17958 956
rect -4480 686 -2600 716
rect -6006 560 -1092 686
rect -6006 -384 -5825 560
rect -5121 -384 -1092 560
rect -6006 -518 -1092 -384
rect 6722 -1734 11058 -1720
rect 5596 -1802 11058 -1734
rect 4386 -1873 5472 -1814
rect 4386 -2075 5030 -1873
rect 4386 -2154 4440 -2075
rect 4396 -2379 4440 -2154
rect 4744 -2097 5030 -2075
rect 5414 -2097 5472 -1873
rect 4744 -2154 5472 -2097
rect 5596 -1895 10810 -1802
rect 4744 -2379 4802 -2154
rect 5596 -2199 6133 -1895
rect 6837 -2199 10810 -1895
rect 5596 -2266 10810 -2199
rect 11034 -2266 11058 -1802
rect 35562 -2042 36656 -2020
rect 5596 -2316 11058 -2266
rect 6722 -2328 11058 -2316
rect 35560 -2054 36656 -2042
rect 38234 -2054 39992 -2020
rect 35560 -2109 39992 -2054
rect 4396 -2514 4802 -2379
rect 35560 -2413 35598 -2109
rect 36222 -2117 39992 -2109
rect 36222 -2413 39125 -2117
rect 35560 -2421 39125 -2413
rect 39909 -2421 39992 -2117
rect 35560 -2488 39992 -2421
rect 35560 -2508 36264 -2488
rect 35576 -2647 36518 -2600
rect 35576 -2791 35697 -2647
rect 36401 -2791 36518 -2647
rect 35576 -2832 36518 -2791
rect -17064 -10702 -8838 -10610
rect -17064 -11406 -9777 -10702
rect -8993 -11406 -8838 -10702
rect -17064 -11570 -8838 -11406
rect -14866 -18164 -13816 -18086
rect -14866 -18720 -14624 -18164
rect -14068 -18720 -13816 -18164
rect -14866 -18812 -13816 -18720
rect 35580 -20279 36510 -20240
rect 35580 -20423 35676 -20279
rect 36460 -20423 36510 -20279
rect 35580 -20466 36510 -20423
rect 94 -21712 490 -21646
rect -2030 -21814 -918 -21810
rect -2030 -22730 -916 -21814
rect -682 -22038 -200 -21804
rect -682 -22662 -597 -22038
rect -293 -22662 -200 -22038
rect 94 -22096 172 -21712
rect 396 -22096 490 -21712
rect 2000 -21693 3122 -21604
rect 2000 -21917 2092 -21693
rect 3036 -21917 3122 -21693
rect 4076 -21674 4296 -21608
rect 2000 -22006 3122 -21917
rect 3254 -21873 3992 -21728
rect 94 -22200 490 -22096
rect 3254 -22382 3359 -21873
rect -2030 -23074 -918 -22730
rect -682 -22782 -200 -22662
rect 3222 -22497 3359 -22382
rect 3903 -22382 3992 -21873
rect 4076 -22298 4117 -21674
rect 4261 -22298 4296 -21674
rect 4076 -22364 4296 -22298
rect 4428 -21772 4626 -21694
rect 4428 -22316 4457 -21772
rect 4601 -21894 4626 -21772
rect 4601 -21987 10228 -21894
rect 4601 -22291 9670 -21987
rect 10134 -22291 10228 -21987
rect 4601 -22316 10228 -22291
rect 3903 -22497 4000 -22382
rect 3222 -22682 4000 -22497
rect -2030 -23858 -1892 -23074
rect -1028 -23858 -918 -23074
rect -2030 -23988 -918 -23858
rect 4084 -24120 4272 -22364
rect 4428 -22404 10228 -22316
rect 4428 -22406 4626 -22404
rect 4084 -24319 5492 -24120
rect 4084 -24555 4377 -24319
rect 4613 -24555 4697 -24319
rect 4933 -24555 5017 -24319
rect 5253 -24555 5492 -24319
rect 4084 -24800 5492 -24555
rect -5992 -24954 -3370 -24940
rect 15082 -24954 39970 -24812
rect -5992 -24969 39970 -24954
rect -5992 -25025 39169 -24969
rect -5992 -25122 3381 -25025
rect -5992 -25906 -5863 -25122
rect -5079 -25889 3381 -25122
rect 3925 -25593 39169 -25025
rect 39793 -25593 39970 -24969
rect 3925 -25889 39970 -25593
rect -5079 -25906 39970 -25889
rect -5992 -25984 39970 -25906
rect -5992 -26000 -3370 -25984
rect 15082 -26070 39970 -25984
rect 11522 -26986 42060 -26922
rect -8000 -27026 42060 -26986
rect -61978 -27151 -53122 -27026
rect -61978 -27855 -60015 -27151
rect -59151 -27855 -53122 -27151
rect -61978 -27986 -53122 -27855
rect -17630 -27054 42060 -27026
rect -17630 -27117 41059 -27054
rect -17630 -27120 2131 -27117
rect -17630 -27904 -7903 -27120
rect -7119 -27901 2131 -27120
rect 2915 -27838 41059 -27117
rect 41763 -27838 42060 -27054
rect 2915 -27901 42060 -27838
rect -7119 -27904 42060 -27901
rect -17630 -27986 42060 -27904
rect -8000 -28014 42060 -27986
rect 11522 -28096 42060 -28014
rect -61946 -29012 12014 -29002
rect -61946 -29124 44086 -29012
rect -61946 -29134 -810 -29124
rect -61946 -29165 -9761 -29134
rect -61946 -29869 -61789 -29165
rect -60925 -29869 -9761 -29165
rect -61946 -29918 -9761 -29869
rect -8977 -29828 -810 -29134
rect -186 -29151 44086 -29124
rect -186 -29828 43199 -29151
rect -8977 -29855 43199 -29828
rect 43823 -29855 44086 -29151
rect -8977 -29918 44086 -29855
rect -61946 -29970 44086 -29918
rect -57840 -30030 44086 -29970
rect 11820 -30036 44086 -30030
<< via4 >>
rect -14624 -18720 -14068 -18164
rect 4377 -24555 4613 -24319
rect 4697 -24555 4933 -24319
rect 5017 -24555 5253 -24319
<< metal5 >>
rect -14866 -18090 -13816 -18086
rect -14866 -18101 -13784 -18090
rect -14866 -18164 -13777 -18101
rect -14866 -18720 -14624 -18164
rect -14068 -18720 -13777 -18164
rect -14866 -18812 -13777 -18720
rect -14834 -18816 -13777 -18812
rect -14471 -24110 -13777 -18816
rect -14471 -24120 4468 -24110
rect -14471 -24319 5492 -24120
rect -14471 -24555 4377 -24319
rect 4613 -24555 4697 -24319
rect 4933 -24555 5017 -24319
rect 5253 -24555 5492 -24319
rect -14471 -24800 5492 -24555
rect -14471 -24804 4468 -24800
use comparator_top  comparator_top_0
timestamp 1686560383
transform 0 -1 8512 1 0 -982
box -7692 -1888 17759 11948
use dac_3v_8bit  dac_3v_8bit_0
timestamp 1686560383
transform 0 -1 35467 -1 0 4301
box -609 -200 25939 24519
use sample_and_hold  sample_and_hold_0
timestamp 1686560383
transform 0 -1 9273 1 0 -21896
box -2224 -1473 19523 12471
use sbamuxm4  sbamuxm4_0
timestamp 1686560383
transform 1 0 -56320 0 1 -10136
box -2839 -17900 44280 24019
<< labels >>
flabel metal4 s -1602 -22484 -1408 -22266 0 FreeSans 14895 0 0 0 vss
port 1 nsew
flabel metal4 s -512 -22482 -348 -22288 0 FreeSans 14895 0 0 0 dvdd
port 2 nsew
flabel metal4 s 232 -22088 298 -22014 0 FreeSans 14895 0 0 0 hold
port 3 nsew
flabel metal4 s 2304 -21882 2436 -21814 0 FreeSans 14895 0 0 0 dvss
port 4 nsew
flabel metal4 s 3504 -22342 3730 -22184 0 FreeSans 14895 0 0 0 vdd
port 5 nsew
flabel metal4 s 4520 -22172 4536 -22040 0 FreeSans 14895 0 0 0 ena
port 6 nsew
flabel metal4 s 4336 11096 4370 11106 0 FreeSans 7627 0 0 0 cmp
port 7 nsew
flabel metal3 s 10792 -10272 10940 -9766 0 FreeSans 6102 0 0 0 dac_out
port 8 nsew
flabel metal4 s 35954 -2762 36128 -2684 0 FreeSans 6102 0 0 0 vhigh
port 9 nsew
flabel metal4 s 35704 -20398 36106 -20338 0 FreeSans 6102 0 0 0 vlow
port 10 nsew
flabel metal4 s 34642 4632 34798 4768 0 FreeSans 6102 0 0 0 b0
port 11 nsew
flabel metal4 s 33010 4678 33166 4814 0 FreeSans 6102 0 0 0 b1
port 12 nsew
flabel metal4 s 31444 4680 31600 4816 0 FreeSans 6102 0 0 0 b2
port 13 nsew
flabel metal4 s 29748 4624 29904 4760 0 FreeSans 6102 0 0 0 b3
port 14 nsew
flabel metal4 s 28216 4698 28372 4834 0 FreeSans 6102 0 0 0 b4
port 15 nsew
flabel metal4 s 26548 4658 26704 4794 0 FreeSans 6102 0 0 0 b5
port 16 nsew
flabel metal4 s 24836 4656 24992 4792 0 FreeSans 6102 0 0 0 b6
port 17 nsew
flabel metal4 s 23182 4634 23338 4770 0 FreeSans 6102 0 0 0 b7
port 18 nsew
flabel metal3 s -56272 -12132 -56244 -12110 0 FreeSans 1562 0 0 0 inp[0]
port 19 nsew
flabel metal3 s -56258 -12528 -56230 -12506 0 FreeSans 1562 0 0 0 inp[1]
port 20 nsew
flabel metal3 s -56224 -12880 -56196 -12858 0 FreeSans 1562 0 0 0 inp[2]
port 21 nsew
flabel metal3 s -56248 -13268 -56220 -13246 0 FreeSans 1562 0 0 0 inp[3]
port 22 nsew
flabel metal3 s -56412 -25282 -56384 -25260 0 FreeSans 1562 0 0 0 inp[4]
port 23 nsew
flabel metal3 s -56382 -25694 -56354 -25672 0 FreeSans 1562 0 0 0 inp[5]
port 24 nsew
flabel metal3 s -56402 -26066 -56374 -26044 0 FreeSans 1562 0 0 0 inp[6]
port 25 nsew
flabel metal3 s -56394 -26442 -56366 -26420 0 FreeSans 1562 0 0 0 inp[7]
port 26 nsew
flabel metal3 s -56658 -16612 -56612 -16558 0 FreeSans 1250 0 0 0 in[0]
port 27 nsew
flabel metal3 s -56550 -19330 -56514 -19298 0 FreeSans 1250 0 0 0 in[1]
port 28 nsew
flabel metal3 s -56564 -21890 -56510 -21854 0 FreeSans 1250 0 0 0 in[2]
port 29 nsew
<< end >>
