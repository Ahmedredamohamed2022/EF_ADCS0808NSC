* NGSPICE file created from EF_ADCS0808NSCM.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_g5v0d10v5_U62SY6 a_n187_n64# w_n387_n362# a_129_n64# a_29_n161#
+ a_n129_n161# a_n29_n64#
X0 a_129_n64# a_29_n161# a_n29_n64# w_n387_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1 a_n29_n64# a_n129_n161# a_n187_n64# w_n387_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EJGQFX a_129_n200# a_29_n288# a_n129_n288# a_n321_n422#
+ a_n29_n200# a_n187_n200#
X0 a_129_n200# a_29_n288# a_n29_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1 a_n29_n200# a_n129_n288# a_n187_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U6NWY6 a_n108_n64# a_50_n64# a_n50_n161# w_n308_n362#
X0 a_50_n64# a_n50_n161# a_n108_n64# w_n308_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8 a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ a_n147_n147# a_n45_n45#
D0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5
.ends

.subckt balanced_switch hold out in vdd vss
Xsky130_fd_pr__pfet_g5v0d10v5_U62SY6_0 holdp vdd holdp holdb holdb vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM1 out holdb holdb vss in out sky130_fd_pr__nfet_g5v0d10v5_EJGQFX
Xsky130_fd_pr__pfet_g5v0d10v5_U6NWY6_0 in in holdb vdd sky130_fd_pr__pfet_g5v0d10v5_U6NWY6
XXM3 in vss in holdp sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
XXM4 out vdd out holdp holdp in sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM5 out vss out holdp sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
XXM6 out out holdb vdd sky130_fd_pr__pfet_g5v0d10v5_U6NWY6
XXM7 holdb vdd holdb hold hold vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM8 holdb vss vss hold sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
XXD1 vss hold sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
XXM10 holdp vss vss holdb sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EJGQJV a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_D7NTZ8 a_n194_2500# a_442_n2932# a_n512_n2932#
+ a_n512_2500# a_n642_n3062# a_124_n2932# a_124_2500# a_442_2500# a_n194_n2932#
X0 a_n194_n2932# a_n194_2500# a_n642_n3062# sky130_fd_pr__res_xhigh_po w=350000u l=2.5e+07u
X1 a_n512_n2932# a_n512_2500# a_n642_n3062# sky130_fd_pr__res_xhigh_po w=350000u l=2.5e+07u
X2 a_442_n2932# a_442_2500# a_n642_n3062# sky130_fd_pr__res_xhigh_po w=350000u l=2.5e+07u
X3 a_124_n2932# a_124_2500# a_n642_n3062# sky130_fd_pr__res_xhigh_po w=350000u l=2.5e+07u
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_EJGQJV a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_03v3_nvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_L93GHW a_n162_n162# a_n60_n60#
D0 a_n162_n162# a_n60_n60# sky130_fd_pr__diode_pw2nd_05v5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT a_n761_n197# a_503_n1069# a_2815_336#
+ a_n129_675# a_1077_336# a_1293_n197# a_n445_n1069# a_n2715_336# a_n977_336# a_2715_n633#
+ a_1709_n100# a_1393_772# a_n2341_239# a_n2973_n633# a_3031_n633# a_n1293_772# a_n2341_n197#
+ a_2025_n100# a_n919_n1069# a_2873_239# a_1925_239# a_1135_n1069# a_n1551_n1069#
+ a_1925_n633# a_1609_n1069# a_1077_n972# a_n1551_n197# a_2241_n633# a_3131_772# a_1235_n100#
+ a_n3031_772# a_n345_772# a_129_336# a_n2715_n536# a_345_n1069# a_445_772# a_n287_n1069#
+ a_n2657_675# a_2241_675# a_n3031_n536# a_2715_n197# a_n1709_675# a_187_239# a_761_n100#
+ a_819_n1069# a_1451_n633# a_2499_n972# a_n2973_n197# a_3031_n197# a_2657_n100# a_n661_n536#
+ a_n1393_n1069# a_287_n536# a_n1925_n536# w_n3389_n1269# a_n2241_n536# a_n1867_n1069#
+ a_1925_n197# a_603_n972# a_2657_336# a_2873_n633# a_n2557_336# a_1709_336# a_2241_n197#
+ a_1867_n100# a_n1609_336# a_n761_n1069# a_2973_772# a_n2183_239# a_n2873_772# a_2183_n100#
+ a_187_n1069# a_n1925_772# a_n1235_239# a_1767_239# a_n1451_n536# a_n1551_675# a_n29_n100#
+ a_1451_n1069# a_1451_n197# a_1709_n972# a_1925_n1069# a_1393_n100# a_2025_n972#
+ a_2025_772# a_n187_772# a_n29_336# a_n2873_n536# a_287_772# a_n603_675# a_1551_336#
+ a_661_n1069# a_n2499_675# a_2083_675# a_n1451_336# a_2873_n197# a_1135_675# a_819_239#
+ a_1235_n972# a_919_n536# a_1293_n1069# a_n187_n100# a_761_n972# a_2499_336# a_1767_n1069#
+ a_n503_336# a_n2399_336# a_2657_n972# a_2815_n100# a_603_336# a_1867_772# a_n2815_239#
+ a_n1077_239# a_n1767_772# a_3131_n100# a_445_n536# a_n1393_675# a_661_239# a_1867_n972#
+ a_977_n1069# a_2183_n972# a_n3189_n100# a_2341_n100# a_n819_772# a_n129_239# a_n2025_n1069#
+ a_n29_n972# a_n3131_675# a_n445_675# a_1393_336# a_919_772# a_n1293_336# a_2715_675#
+ a_1393_n972# a_n2399_n100# a_1551_n100# a_977_675# a_n819_n100# a_1077_n536# a_3131_336#
+ a_n3031_336# a_n345_336# a_2973_n100# a_29_n633# a_n661_772# a_445_336# a_n2657_239#
+ a_2241_239# a_n1709_239# a_761_772# a_n187_n972# a_2499_n536# a_n2973_675# a_n345_n100#
+ a_n129_n633# a_n1609_n100# a_2815_n972# a_3131_n972# a_603_n536# a_n2341_n1069#
+ a_2973_336# a_187_n633# a_n287_675# a_n2025_675# a_n2873_336# a_2557_675# a_n1925_336#
+ a_1609_675# a_29_n197# a_n3189_n972# a_n2815_n1069# a_n1135_n100# a_2341_n972# a_n1551_239#
+ a_1709_n536# a_n977_n100# a_n129_n197# a_2025_n536# a_2025_336# a_n2399_n972# a_n187_336#
+ a_1551_n972# a_n2557_n100# a_2341_772# a_29_675# a_n2241_772# a_n603_239# a_287_336#
+ a_n2499_239# a_2083_239# a_n2183_n1069# a_n819_n972# a_1135_239# a_187_n197# a_1235_n536#
+ a_n1867_675# a_1451_675# a_n287_n633# a_n2657_n1069# a_n1767_n100# a_2973_n972#
+ a_n2083_n100# a_761_n536# a_n3189_772# a_819_n633# a_n345_n972# a_2657_n536# a_n503_n100#
+ a_2241_n1069# a_n919_675# a_n1609_n972# a_1867_336# a_2399_675# a_n1767_336# a_129_n100#
+ a_n1293_n100# a_n1393_239# a_n1077_n633# a_2715_n1069# a_503_675# a_1867_n536# a_n2499_n1069#
+ a_345_n633# a_2183_n536# a_n287_n197# a_n1135_n972# a_n819_336# a_2183_772# a_n3131_239#
+ a_n2499_n633# a_n29_n536# a_n2083_772# a_1235_772# a_n445_239# a_n1135_772# a_919_336#
+ a_n977_n972# a_2715_239# a_819_n197# a_n761_675# a_2083_n1069# a_1393_n536# a_n919_n633#
+ a_1293_675# a_977_239# a_n2557_n972# a_2557_n1069# a_n2973_n1069# a_n2715_n100#
+ a_n1077_n197# a_n3031_n100# a_977_n633# a_345_n197# a_n661_n100# a_3031_675# a_n661_336#
+ a_n1767_n972# a_n445_n633# a_287_n100# a_n1925_n100# a_n2083_n972# a_761_336# a_n2499_n197#
+ a_n1709_n633# a_n2973_239# a_n187_n536# a_n2241_n100# a_29_n1069# a_345_675# a_n2025_n633#
+ a_n919_n197# a_n503_n972# a_2815_n536# a_2399_n1069# a_129_n972# a_3131_n536# a_n1293_n972#
+ a_2399_n633# a_n1451_n100# a_n1235_n633# a_2815_772# a_n977_772# a_1077_772# a_n2025_239#
+ a_n287_239# a_n2715_772# a_977_n197# a_2557_239# a_n2341_675# a_1609_239# a_n3189_n536#
+ a_503_n633# a_2341_n536# a_2873_675# a_n445_n197# a_1925_675# a_n1709_n197# a_n2873_n100#
+ a_n2657_n633# a_2873_n1069# a_n2025_n197# a_n2399_n536# a_1551_n536# a_29_239# a_2341_336#
+ a_129_772# a_919_n100# a_n2241_336# a_2399_n197# a_1609_n633# a_n2715_n972# a_n819_n536#
+ a_n1867_n633# a_n1235_n197# a_n3031_n972# a_187_675# a_n1867_239# a_n2183_n633#
+ a_1451_239# a_n661_n972# a_2973_n536# a_503_n197# a_287_n972# a_n3131_n1069# a_n1925_n972#
+ a_n603_n633# a_445_n100# a_n3189_336# a_1135_n633# a_n2241_n972# a_n2657_n197# a_n345_n536#
+ a_n1393_n633# a_2657_772# a_n2557_772# a_1709_772# a_n919_239# a_n1609_n536# a_n1609_772#
+ a_2399_239# a_n2183_675# a_661_n633# a_n1235_675# a_1609_n197# a_503_239# a_1767_675#
+ a_n1451_n972# a_n1867_n197# a_2557_n633# a_n2183_n197# a_n1135_n536# a_n129_n1069#
+ a_2183_336# a_n603_n197# a_n2083_336# a_1767_n633# a_n29_772# a_1235_336# a_1135_n197#
+ a_n2873_n972# a_n1135_336# a_n977_n536# a_n1393_n197# a_2083_n633# a_1551_772# a_n761_239#
+ a_1077_n100# a_n2815_n633# a_n1451_772# a_n1235_n1069# a_819_675# a_1293_239# a_n3131_n633#
+ a_n2557_n536# a_661_n197# a_919_n972# a_n1709_n1069# a_n761_n633# a_2557_n197# a_3031_n1069#
+ a_1293_n633# a_2499_n100# a_n603_n1069# a_n503_772# a_2499_772# a_n2341_n633# a_3031_239#
+ a_n2399_772# a_n1767_n536# a_603_772# a_n2083_n536# a_n2815_675# a_1767_n197# a_445_n972#
+ a_n1077_675# a_345_239# a_603_n100# a_2083_n197# a_661_675# a_n2815_n197# a_n1077_n1069#
+ a_n503_n536# a_n1551_n633# a_n3131_n197# a_129_n536# a_n1293_n536#
X0 a_n2557_772# a_n2657_675# a_n2715_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1 a_287_n100# a_187_n197# a_129_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2 a_1709_n100# a_1609_n197# a_1551_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3 a_1077_772# a_977_675# a_919_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4 a_n2083_772# a_n2183_675# a_n2241_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X5 a_1235_n100# a_1135_n197# a_1077_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X6 a_2025_772# a_1925_675# a_1867_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X7 a_n1925_336# a_n2025_239# a_n2083_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X8 a_919_336# a_819_239# a_761_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X9 a_1551_772# a_1451_675# a_1393_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X10 a_445_336# a_345_239# a_287_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X11 a_n977_n972# a_n1077_n1069# a_n1135_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X12 a_919_n100# a_819_n197# a_761_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X13 a_n1925_n100# a_n2025_n197# a_n2083_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X14 a_445_n100# a_345_n197# a_287_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X15 a_n2715_772# a_n2815_675# a_n2873_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X16 a_1077_n972# a_977_n1069# a_919_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X17 a_n2241_772# a_n2341_675# a_n2399_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X18 a_n503_n972# a_n603_n1069# a_n661_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X19 a_3131_336# a_3031_239# a_2973_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X20 a_2657_n972# a_2557_n1069# a_2499_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X21 a_1235_n536# a_1135_n633# a_1077_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X22 a_n1135_n536# a_n1235_n633# a_n1293_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X23 a_761_772# a_661_675# a_603_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X24 a_n2557_n972# a_n2657_n1069# a_n2715_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X25 a_603_336# a_503_239# a_445_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X26 a_3131_n100# a_3031_n197# a_2973_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X27 a_603_n100# a_503_n197# a_445_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X28 a_2815_n536# a_2715_n633# a_2657_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X29 a_n2715_n536# a_n2815_n633# a_n2873_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X30 a_287_772# a_187_675# a_129_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X31 a_1709_772# a_1609_675# a_1551_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X32 a_603_n972# a_503_n1069# a_445_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X33 a_n29_n972# a_n129_n1069# a_n187_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X34 a_1235_772# a_1135_675# a_1077_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X35 a_3131_n536# a_3031_n633# a_2973_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X36 a_n3031_n536# a_n3131_n633# a_n3189_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X37 a_n1925_772# a_n2025_675# a_n2083_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X38 a_919_772# a_819_675# a_761_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X39 a_n1767_336# a_n1867_239# a_n1925_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X40 a_445_772# a_345_675# a_287_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X41 a_n1293_336# a_n1393_239# a_n1451_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X42 a_1867_n536# a_1767_n633# a_1709_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X43 a_n1767_n536# a_n1867_n633# a_n1925_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X44 a_n1767_n100# a_n1867_n197# a_n1925_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X45 a_n1293_n100# a_n1393_n197# a_n1451_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X46 a_2183_n536# a_2083_n633# a_2025_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X47 a_n2083_n536# a_n2183_n633# a_n2241_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X48 a_3131_772# a_3031_675# a_2973_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X49 a_2973_336# a_2873_239# a_2815_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X50 a_1235_n972# a_1135_n1069# a_1077_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X51 a_n1135_n972# a_n1235_n1069# a_n1293_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X52 a_603_772# a_503_675# a_445_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X53 a_n1451_336# a_n1551_239# a_n1609_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X54 a_2973_n100# a_2873_n197# a_2815_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X55 a_2815_n972# a_2715_n1069# a_2657_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X56 a_n2715_n972# a_n2815_n1069# a_n2873_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X57 a_2499_336# a_2399_239# a_2341_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X58 a_n1451_n100# a_n1551_n197# a_n1609_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X59 a_n819_n536# a_n919_n633# a_n977_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X60 a_n977_336# a_n1077_239# a_n1135_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X61 a_3131_n972# a_3031_n1069# a_2973_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X62 a_n3031_n972# a_n3131_n1069# a_n3189_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X63 a_2499_n100# a_2399_n197# a_2341_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X64 a_n661_n536# a_n761_n633# a_n819_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X65 a_n977_n100# a_n1077_n197# a_n1135_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X66 a_n1767_772# a_n1867_675# a_n1925_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X67 a_2657_336# a_2557_239# a_2499_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X68 a_n1609_336# a_n1709_239# a_n1767_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X69 a_1867_n972# a_1767_n1069# a_1709_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X70 a_n1767_n972# a_n1867_n1069# a_n1925_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X71 a_n1293_772# a_n1393_675# a_n1451_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X72 a_2183_336# a_2083_239# a_2025_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X73 a_n1135_336# a_n1235_239# a_n1293_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X74 a_919_n536# a_819_n633# a_761_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X75 a_2657_n100# a_2557_n197# a_2499_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X76 a_n1609_n100# a_n1709_n197# a_n1767_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X77 a_2183_n972# a_2083_n1069# a_2025_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X78 a_2183_n100# a_2083_n197# a_2025_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X79 a_n2083_n972# a_n2183_n1069# a_n2241_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X80 a_2025_n536# a_1925_n633# a_1867_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X81 a_2973_772# a_2873_675# a_2815_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X82 a_n1135_n100# a_n1235_n197# a_n1293_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X83 a_761_n536# a_661_n633# a_603_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X84 a_n187_n536# a_n287_n633# a_n345_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X85 a_2815_336# a_2715_239# a_2657_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X86 a_n1451_772# a_n1551_675# a_n1609_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X87 a_2341_336# a_2241_239# a_2183_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X88 a_2341_n536# a_2241_n633# a_2183_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X89 a_n2241_n536# a_n2341_n633# a_n2399_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X90 a_2815_n100# a_2715_n197# a_2657_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X91 a_2499_772# a_2399_675# a_2341_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X92 a_n661_336# a_n761_239# a_n819_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X93 a_2341_n100# a_2241_n197# a_2183_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X94 a_n3031_336# a_n3131_239# a_n3189_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X95 a_n819_n972# a_n919_n1069# a_n977_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X96 a_n977_772# a_n1077_675# a_n1135_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X97 a_129_336# a_29_239# a_n29_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X98 a_n661_n100# a_n761_n197# a_n819_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X99 a_287_n536# a_187_n633# a_129_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X100 a_n3031_n100# a_n3131_n197# a_n3189_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X101 a_129_n100# a_29_n197# a_n29_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X102 a_n661_n972# a_n761_n1069# a_n819_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X103 a_n187_336# a_n287_239# a_n345_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X104 a_1393_n536# a_1293_n633# a_1235_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X105 a_n1293_n536# a_n1393_n633# a_n1451_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X106 a_2657_772# a_2557_675# a_2499_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X107 a_n1609_772# a_n1709_675# a_n1767_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X108 a_2183_772# a_2083_675# a_2025_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X109 a_n187_n100# a_n287_n197# a_n345_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X110 a_n1135_772# a_n1235_675# a_n1293_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X111 a_919_n972# a_819_n1069# a_761_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X112 a_n819_336# a_n919_239# a_n977_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X113 a_2973_n536# a_2873_n633# a_2815_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X114 a_n2873_n536# a_n2973_n633# a_n3031_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X115 a_2025_n972# a_1925_n1069# a_1867_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X116 a_n345_336# a_n445_239# a_n503_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X117 a_761_n972# a_661_n1069# a_603_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X118 a_n187_n972# a_n287_n1069# a_n345_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X119 a_2815_772# a_2715_675# a_2657_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X120 a_n819_n100# a_n919_n197# a_n977_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X121 a_2341_772# a_2241_675# a_2183_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X122 a_n345_n100# a_n445_n197# a_n503_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X123 a_2341_n972# a_2241_n1069# a_2183_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X124 a_n2241_n972# a_n2341_n1069# a_n2399_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X125 a_n345_n536# a_n445_n633# a_n503_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X126 a_n661_772# a_n761_675# a_n819_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X127 a_2499_n536# a_2399_n633# a_2341_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X128 a_n2399_n536# a_n2499_n633# a_n2557_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X129 a_n3031_772# a_n3131_675# a_n3189_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X130 a_n2873_336# a_n2973_239# a_n3031_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X131 a_n503_336# a_n603_239# a_n661_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X132 a_129_772# a_29_675# a_n29_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X133 a_287_n972# a_187_n1069# a_129_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X134 a_n503_n100# a_n603_n197# a_n661_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X135 a_129_n536# a_29_n633# a_n29_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X136 a_n2873_n100# a_n2973_n197# a_n3031_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X137 a_n187_772# a_n287_675# a_n345_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X138 a_1393_n972# a_1293_n1069# a_1235_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X139 a_n1293_n972# a_n1393_n1069# a_n1451_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X140 a_1709_n536# a_1609_n633# a_1551_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X141 a_n1609_n536# a_n1709_n633# a_n1767_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X142 a_n2399_336# a_n2499_239# a_n2557_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X143 a_n29_336# a_n129_239# a_n187_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X144 a_445_n536# a_345_n633# a_287_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X145 a_n29_n100# a_n129_n197# a_n187_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X146 a_1867_336# a_1767_239# a_1709_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X147 a_n2399_n100# a_n2499_n197# a_n2557_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X148 a_1551_n536# a_1451_n633# a_1393_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X149 a_n1451_n536# a_n1551_n633# a_n1609_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X150 a_n1925_n536# a_n2025_n633# a_n2083_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X151 a_n819_772# a_n919_675# a_n977_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X152 a_2973_n972# a_2873_n1069# a_2815_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X153 a_n2873_n972# a_n2973_n1069# a_n3031_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X154 a_1393_336# a_1293_239# a_1235_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X155 a_n345_772# a_n445_675# a_n503_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X156 a_1867_n100# a_1767_n197# a_1709_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X157 a_n2557_336# a_n2657_239# a_n2715_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X158 a_1393_n100# a_1293_n197# a_1235_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X159 a_1077_336# a_977_239# a_919_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X160 a_n2083_336# a_n2183_239# a_n2241_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X161 a_2025_336# a_1925_239# a_1867_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X162 a_n2557_n100# a_n2657_n197# a_n2715_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X163 a_n345_n972# a_n445_n1069# a_n503_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X164 a_1551_336# a_1451_239# a_1393_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X165 a_n2083_n100# a_n2183_n197# a_n2241_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X166 a_1077_n100# a_977_n197# a_919_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X167 a_2499_n972# a_2399_n1069# a_2341_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X168 a_n977_n536# a_n1077_n633# a_n1135_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X169 a_n2873_772# a_n2973_675# a_n3031_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X170 a_n503_772# a_n603_675# a_n661_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X171 a_n2399_n972# a_n2499_n1069# a_n2557_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X172 a_2025_n100# a_1925_n197# a_1867_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X173 a_n2715_336# a_n2815_239# a_n2873_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X174 a_1077_n536# a_977_n633# a_919_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X175 a_1551_n100# a_1451_n197# a_1393_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X176 a_n2241_336# a_n2341_239# a_n2399_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X177 a_n503_n536# a_n603_n633# a_n661_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X178 a_129_n972# a_29_n1069# a_n29_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X179 a_2657_n536# a_2557_n633# a_2499_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X180 a_761_336# a_661_239# a_603_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X181 a_n2715_n100# a_n2815_n197# a_n2873_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X182 a_n2557_n536# a_n2657_n633# a_n2715_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X183 a_1709_n972# a_1609_n1069# a_1551_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X184 a_n2399_772# a_n2499_675# a_n2557_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X185 a_n29_772# a_n129_675# a_n187_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X186 a_n2241_n100# a_n2341_n197# a_n2399_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X187 a_n1609_n972# a_n1709_n1069# a_n1767_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X188 a_445_n972# a_345_n1069# a_287_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X189 a_761_n100# a_661_n197# a_603_n100# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X190 a_1867_772# a_1767_675# a_1709_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X191 a_1551_n972# a_1451_n1069# a_1393_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X192 a_n1451_n972# a_n1551_n1069# a_n1609_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X193 a_n1925_n972# a_n2025_n1069# a_n2083_n972# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X194 a_287_336# a_187_239# a_129_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X195 a_1709_336# a_1609_239# a_1551_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X196 a_1393_772# a_1293_675# a_1235_772# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X197 a_603_n536# a_503_n633# a_445_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X198 a_n29_n536# a_n129_n633# a_n187_n536# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X199 a_1235_336# a_1135_239# a_1077_336# w_n3389_n1269# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_H7BQ24 a_n287_n188# a_n29_n100# a_n187_n100#
+ a_n345_n100# a_129_n100# a_287_n100# a_n479_n322# a_29_n188# a_n129_n188# a_187_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1 a_n187_n100# a_n287_n188# a_n345_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2 a_n29_n100# a_n129_n188# a_n187_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3 a_287_n100# a_187_n188# a_129_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UC3VEF a_n1077_230# a_n2815_230# a_1709_n100#
+ a_n1077_n606# a_2025_n100# a_661_230# a_345_n606# a_n2715_n518# a_129_318# a_n2499_n606#
+ a_n3031_n518# a_n129_230# a_1235_n100# a_n661_n518# a_n287_n188# a_n919_n606# a_287_n518#
+ a_n1925_n518# a_n2241_n518# a_761_n100# a_2657_n100# a_819_n188# a_2657_318# a_n2557_318#
+ a_977_n606# a_1709_318# a_n1609_318# a_n445_n606# a_n1451_n518# a_n1077_n188# a_n1709_n606#
+ a_2241_230# a_n2657_230# a_1867_n100# a_n2025_n606# a_n1709_230# a_2183_n100# a_345_n188#
+ a_2399_n606# a_n2873_n518# a_n29_n100# a_n2499_n188# a_n29_318# a_n1235_n606# a_1551_318#
+ a_n1451_318# a_1393_n100# a_n919_n188# a_503_n606# a_919_n518# a_n1551_230# a_n2657_n606#
+ a_977_n188# a_2499_318# a_n503_318# a_n2399_318# a_n445_n188# a_603_318# a_1609_n606#
+ a_445_n518# a_n1709_n188# a_n1867_n606# a_n187_n100# a_n603_230# a_n2025_n188# a_2083_230#
+ a_n2499_230# a_2815_n100# a_n2183_n606# a_1135_230# a_3131_n100# a_n603_n606# a_2399_n188#
+ a_1135_n606# a_n1235_n188# a_n1393_n606# a_1393_318# a_n1293_318# a_n3189_n100#
+ a_503_n188# a_2341_n100# a_661_n606# a_2557_n606# a_1077_n518# a_n2657_n188# a_n1393_230#
+ a_3131_318# a_n3031_318# a_1551_n100# a_n2399_n100# a_n345_318# a_1609_n188# a_445_318#
+ a_1767_n606# a_n819_n100# a_n1867_n188# a_2083_n606# a_2499_n518# a_n2183_n188#
+ a_n445_230# a_n3131_230# a_n2815_n606# a_2715_230# a_2973_n100# a_n3131_n606# a_n603_n188#
+ a_977_230# a_n761_n606# a_603_n518# a_1135_n188# a_1293_n606# a_n345_n100# a_n1393_n188#
+ a_n2341_n606# a_n1609_n100# a_2973_318# a_n2873_318# a_661_n188# a_n1925_318# a_2557_n188#
+ a_1709_n518# a_n2973_230# a_n1551_n606# a_2025_n518# a_2025_318# a_n1135_n100# a_n187_318#
+ a_1767_n188# a_287_318# a_2715_n606# a_n977_n100# a_2083_n188# a_n2815_n188# a_n2973_n606#
+ a_1235_n518# a_n287_230# a_n2025_230# a_3031_n606# a_n2557_n100# a_n3131_n188# a_2557_230#
+ a_1609_230# a_761_n518# a_1293_n188# a_n761_n188# a_1925_n606# a_2241_n606# a_2657_n518#
+ a_n2341_n188# a_n1767_n100# a_1867_318# a_n2083_n100# a_n1767_318# a_29_230# a_1451_n606#
+ a_1867_n518# a_n1551_n188# a_2183_n518# a_n503_n100# a_1451_230# a_n1867_230# a_129_n100#
+ a_n1293_n100# a_n29_n518# a_n819_318# a_2715_n188# a_919_318# a_2873_n606# a_3031_n188#
+ a_n2973_n188# a_1393_n518# a_n919_230# a_2399_230# a_1925_n188# a_503_230# a_2241_n188#
+ a_n661_318# a_n2715_n100# a_n187_n518# a_n3031_n100# a_761_318# a_1451_n188# a_2815_n518#
+ a_n661_n100# a_n761_230# a_287_n100# a_n1925_n100# a_1293_230# a_3131_n518# a_n2241_n100#
+ a_2873_n188# a_n3189_n518# a_2341_n518# a_3031_230# a_n1451_n100# a_345_230# a_n2399_n518#
+ a_1551_n518# a_2341_318# a_n2241_318# a_n819_n518# a_n2873_n100# a_919_n100# a_2973_n518#
+ a_n2341_230# a_2873_230# a_1925_230# a_n3189_318# a_n345_n518# a_n3323_n740# a_n1609_n518#
+ a_29_n606# a_445_n100# a_187_230# a_n129_n606# a_n1135_n518# a_2183_318# a_1235_318#
+ a_n2083_318# a_n977_n518# a_n1135_318# a_187_n606# a_n2557_n518# a_n1235_230# a_n2183_230#
+ a_1767_230# a_1077_n100# a_n1767_n518# a_29_n188# a_n2083_n518# a_2499_n100# a_n503_n518#
+ a_n129_n188# a_n287_n606# a_n1293_n518# a_129_n518# a_819_230# a_603_n100# a_2815_318#
+ a_1077_318# a_n977_318# a_n2715_318# a_187_n188# a_819_n606#
X0 a_1709_n518# a_1609_n606# a_1551_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1 a_n1609_n518# a_n1709_n606# a_n1767_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2 a_n2399_318# a_n2499_230# a_n2557_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3 a_n29_318# a_n129_230# a_n187_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4 a_445_n518# a_345_n606# a_287_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X5 a_919_n100# a_819_n188# a_761_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X6 a_n1925_n100# a_n2025_n188# a_n2083_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X7 a_445_n100# a_345_n188# a_287_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X8 a_1551_n518# a_1451_n606# a_1393_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X9 a_n1451_n518# a_n1551_n606# a_n1609_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X10 a_n1925_n518# a_n2025_n606# a_n2083_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X11 a_1867_318# a_1767_230# a_1709_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X12 a_1393_318# a_1293_230# a_1235_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X13 a_n2557_318# a_n2657_230# a_n2715_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X14 a_3131_n100# a_3031_n188# a_2973_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X15 a_1077_318# a_977_230# a_919_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X16 a_n2083_318# a_n2183_230# a_n2241_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X17 a_603_n100# a_503_n188# a_445_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X18 a_2025_318# a_1925_230# a_1867_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X19 a_1551_318# a_1451_230# a_1393_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X20 a_n977_n518# a_n1077_n606# a_n1135_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X21 a_n2715_318# a_n2815_230# a_n2873_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X22 a_1077_n518# a_977_n606# a_919_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X23 a_n2241_318# a_n2341_230# a_n2399_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X24 a_n503_n518# a_n603_n606# a_n661_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X25 a_2657_n518# a_2557_n606# a_2499_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X26 a_n2557_n518# a_n2657_n606# a_n2715_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X27 a_761_318# a_661_230# a_603_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X28 a_n1767_n100# a_n1867_n188# a_n1925_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X29 a_n1293_n100# a_n1393_n188# a_n1451_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X30 a_287_318# a_187_230# a_129_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X31 a_1709_318# a_1609_230# a_1551_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X32 a_603_n518# a_503_n606# a_445_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X33 a_n29_n518# a_n129_n606# a_n187_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X34 a_1235_318# a_1135_230# a_1077_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X35 a_2973_n100# a_2873_n188# a_2815_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X36 a_n1925_318# a_n2025_230# a_n2083_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X37 a_n1451_n100# a_n1551_n188# a_n1609_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X38 a_919_318# a_819_230# a_761_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X39 a_445_318# a_345_230# a_287_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X40 a_2499_n100# a_2399_n188# a_2341_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X41 a_1235_n518# a_1135_n606# a_1077_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X42 a_n977_n100# a_n1077_n188# a_n1135_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X43 a_n1135_n518# a_n1235_n606# a_n1293_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X44 a_3131_318# a_3031_230# a_2973_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X45 a_603_318# a_503_230# a_445_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X46 a_2657_n100# a_2557_n188# a_2499_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X47 a_2815_n518# a_2715_n606# a_2657_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X48 a_n2715_n518# a_n2815_n606# a_n2873_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X49 a_n1609_n100# a_n1709_n188# a_n1767_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X50 a_2183_n100# a_2083_n188# a_2025_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X51 a_n1135_n100# a_n1235_n188# a_n1293_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X52 a_3131_n518# a_3031_n606# a_2973_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X53 a_n3031_n518# a_n3131_n606# a_n3189_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X54 a_2815_n100# a_2715_n188# a_2657_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X55 a_n1767_318# a_n1867_230# a_n1925_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X56 a_1867_n518# a_1767_n606# a_1709_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X57 a_2341_n100# a_2241_n188# a_2183_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X58 a_n1293_318# a_n1393_230# a_n1451_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X59 a_n1767_n518# a_n1867_n606# a_n1925_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X60 a_n661_n100# a_n761_n188# a_n819_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X61 a_2183_n518# a_2083_n606# a_2025_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X62 a_n2083_n518# a_n2183_n606# a_n2241_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X63 a_n3031_n100# a_n3131_n188# a_n3189_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X64 a_129_n100# a_29_n188# a_n29_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X65 a_2973_318# a_2873_230# a_2815_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X66 a_n1451_318# a_n1551_230# a_n1609_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X67 a_n187_n100# a_n287_n188# a_n345_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X68 a_2499_318# a_2399_230# a_2341_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X69 a_n819_n518# a_n919_n606# a_n977_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X70 a_n977_318# a_n1077_230# a_n1135_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X71 a_n819_n100# a_n919_n188# a_n977_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X72 a_n345_n100# a_n445_n188# a_n503_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X73 a_n661_n518# a_n761_n606# a_n819_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X74 a_2657_318# a_2557_230# a_2499_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X75 a_n1609_318# a_n1709_230# a_n1767_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X76 a_2183_318# a_2083_230# a_2025_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X77 a_n1135_318# a_n1235_230# a_n1293_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X78 a_919_n518# a_819_n606# a_761_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X79 a_n503_n100# a_n603_n188# a_n661_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X80 a_n2873_n100# a_n2973_n188# a_n3031_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X81 a_2025_n518# a_1925_n606# a_1867_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X82 a_761_n518# a_661_n606# a_603_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X83 a_n187_n518# a_n287_n606# a_n345_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X84 a_2815_318# a_2715_230# a_2657_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X85 a_2341_n518# a_2241_n606# a_2183_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X86 a_2341_318# a_2241_230# a_2183_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X87 a_n2241_n518# a_n2341_n606# a_n2399_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X88 a_n29_n100# a_n129_n188# a_n187_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X89 a_n2399_n100# a_n2499_n188# a_n2557_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X90 a_n661_318# a_n761_230# a_n819_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X91 a_n3031_318# a_n3131_230# a_n3189_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X92 a_1867_n100# a_1767_n188# a_1709_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X93 a_129_318# a_29_230# a_n29_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X94 a_287_n518# a_187_n606# a_129_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X95 a_1393_n100# a_1293_n188# a_1235_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X96 a_n187_318# a_n287_230# a_n345_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X97 a_1393_n518# a_1293_n606# a_1235_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X98 a_n2557_n100# a_n2657_n188# a_n2715_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X99 a_n1293_n518# a_n1393_n606# a_n1451_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X100 a_1077_n100# a_977_n188# a_919_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X101 a_n2083_n100# a_n2183_n188# a_n2241_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X102 a_2025_n100# a_1925_n188# a_1867_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X103 a_1551_n100# a_1451_n188# a_1393_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X104 a_2973_n518# a_2873_n606# a_2815_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X105 a_n819_318# a_n919_230# a_n977_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X106 a_n2873_n518# a_n2973_n606# a_n3031_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X107 a_n345_318# a_n445_230# a_n503_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X108 a_n2715_n100# a_n2815_n188# a_n2873_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X109 a_n2241_n100# a_n2341_n188# a_n2399_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X110 a_761_n100# a_661_n188# a_603_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X111 a_n345_n518# a_n445_n606# a_n503_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X112 a_2499_n518# a_2399_n606# a_2341_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X113 a_n2399_n518# a_n2499_n606# a_n2557_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X114 a_n2873_318# a_n2973_230# a_n3031_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X115 a_n503_318# a_n603_230# a_n661_318# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X116 a_1709_n100# a_1609_n188# a_1551_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X117 a_287_n100# a_187_n188# a_129_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X118 a_129_n518# a_29_n606# a_n29_n518# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X119 a_1235_n100# a_1135_n188# a_1077_n100# a_n3323_n740# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
.ends

.subckt follower_amp vdd in out ena vss
XXM25 vdd pbias pbias vdd sky130_fd_pr__pfet_g5v0d10v5_U6NWY6
XXM26 vcomp vdd vcomp pbias pbias vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM27 m1_n523_n317# vdd m1_n523_n317# out out vcomp sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM28 ndrv vdd ndrv in in vcomp sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XM13 m1_1604_n2434# vss nbias ena sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
XM24 vss vss pbias nbias sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
XXM29 ndrv vss vss m1_n523_n317# sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
Xsky130_fd_pr__res_xhigh_po_0p35_D7NTZ8_0 m1_1621_n3043# m1_n3792_n3361# m1_n3792_n2735#
+ m1_1604_n2434# vss m1_n3792_n3361# m1_1621_n3043# vdd m1_n3792_n2735# sky130_fd_pr__res_xhigh_po_0p35_D7NTZ8
XXM1 vcomn1 vss m1_n1946_423# out sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
XXM2 vcomn1 vss pdrv1 in sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
XXM3 pdrv2 vdd pdrv2 m1_n3113_423# m1_n3113_423# vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM4 pdrv1 vdd pdrv1 m1_n1946_423# m1_n1946_423# vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM5 m1_n1946_423# vdd m1_n1946_423# m1_n1946_423# m1_n1946_423# vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM6 m1_n3113_423# vdd m1_n3113_423# m1_n3113_423# m1_n3113_423# vdd sky130_fd_pr__pfet_g5v0d10v5_U62SY6
XXM7 vss vss vcomn2 nbias sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
XXM9 vss vss vcomn1 nbias sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
XXM8 vcomn2 vss m1_n3113_423# out sky130_fd_pr__nfet_03v3_nvt_EJGQJV
Xsky130_fd_pr__nfet_03v3_nvt_EJGQJV_0 vcomn2 vss pdrv2 in sky130_fd_pr__nfet_03v3_nvt_EJGQJV
Xsky130_fd_pr__diode_pw2nd_05v5_L93GHW_0 vss ena sky130_fd_pr__diode_pw2nd_05v5_L93GHW
Xsky130_fd_pr__diode_pw2nd_05v5_L93GHW_1 vss in sky130_fd_pr__diode_pw2nd_05v5_L93GHW
Xsky130_fd_pr__pfet_g5v0d10v5_AQ2AJT_0 pdrv1 pdrv1 out pdrv1 vdd pdrv1 pdrv1 vdd out
+ pdrv1 vdd vdd pdrv1 pdrv1 pdrv1 out pdrv1 vdd pdrv1 pdrv1 pdrv1 pdrv1 pdrv1 pdrv1
+ pdrv1 vdd pdrv1 pdrv1 out out vdd out vdd vdd pdrv1 vdd pdrv1 pdrv1 pdrv1 vdd pdrv1
+ pdrv1 pdrv1 vdd pdrv1 pdrv1 out pdrv1 pdrv1 vdd out pdrv1 out out vdd out pdrv1
+ pdrv1 out vdd pdrv1 out vdd pdrv1 out out pdrv1 vdd pdrv1 out out pdrv1 out pdrv1
+ pdrv1 vdd pdrv1 out pdrv1 pdrv1 vdd pdrv1 vdd vdd vdd vdd out out out pdrv1 out
+ pdrv1 pdrv1 pdrv1 vdd pdrv1 pdrv1 pdrv1 out out pdrv1 vdd vdd out pdrv1 vdd vdd
+ vdd out out out pdrv1 pdrv1 vdd out vdd pdrv1 pdrv1 out pdrv1 out out vdd vdd pdrv1
+ pdrv1 out pdrv1 pdrv1 vdd out out pdrv1 vdd vdd out pdrv1 vdd vdd out vdd out vdd
+ pdrv1 out vdd pdrv1 pdrv1 pdrv1 vdd vdd out pdrv1 out pdrv1 out out out out pdrv1
+ vdd pdrv1 pdrv1 pdrv1 out pdrv1 out pdrv1 pdrv1 out pdrv1 vdd vdd pdrv1 vdd out
+ pdrv1 vdd vdd vdd vdd out out vdd pdrv1 out pdrv1 out pdrv1 pdrv1 pdrv1 vdd pdrv1
+ pdrv1 out pdrv1 pdrv1 pdrv1 pdrv1 vdd vdd vdd vdd out pdrv1 out vdd vdd pdrv1 pdrv1
+ out out pdrv1 vdd vdd out pdrv1 pdrv1 pdrv1 pdrv1 out pdrv1 pdrv1 out pdrv1 vdd
+ vdd out pdrv1 pdrv1 out vdd out pdrv1 vdd out out pdrv1 pdrv1 pdrv1 pdrv1 vdd pdrv1
+ pdrv1 pdrv1 out pdrv1 pdrv1 vdd pdrv1 vdd pdrv1 pdrv1 out pdrv1 out vdd pdrv1 out
+ out vdd vdd pdrv1 pdrv1 pdrv1 vdd out pdrv1 pdrv1 pdrv1 pdrv1 vdd out pdrv1 vdd
+ out out pdrv1 vdd pdrv1 out out vdd pdrv1 pdrv1 vdd pdrv1 pdrv1 pdrv1 pdrv1 out
+ pdrv1 vdd pdrv1 pdrv1 pdrv1 pdrv1 out pdrv1 pdrv1 pdrv1 vdd out pdrv1 vdd vdd out
+ out pdrv1 pdrv1 vdd vdd pdrv1 pdrv1 vdd pdrv1 pdrv1 pdrv1 pdrv1 out vdd pdrv1 out
+ pdrv1 out pdrv1 vdd out pdrv1 out pdrv1 out pdrv1 vdd out vdd pdrv1 out out pdrv1
+ pdrv1 pdrv1 pdrv1 pdrv1 pdrv1 pdrv1 vdd pdrv1 pdrv1 pdrv1 vdd pdrv1 out pdrv1 vdd
+ pdrv1 out out pdrv1 out vdd out pdrv1 pdrv1 out pdrv1 vdd pdrv1 vdd pdrv1 pdrv1
+ pdrv1 pdrv1 out pdrv1 out pdrv1 pdrv1 pdrv1 pdrv1 pdrv1 out pdrv1 vdd out pdrv1
+ pdrv1 vdd vdd out vdd pdrv1 pdrv1 vdd pdrv1 pdrv1 out pdrv1 pdrv1 pdrv1 pdrv1 vdd
+ pdrv1 pdrv1 vdd out sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT
Xsky130_fd_pr__pfet_g5v0d10v5_AQ2AJT_1 pdrv2 pdrv2 out pdrv2 vdd pdrv2 pdrv2 vdd out
+ pdrv2 vdd vdd pdrv2 pdrv2 pdrv2 out pdrv2 vdd pdrv2 pdrv2 pdrv2 pdrv2 pdrv2 pdrv2
+ pdrv2 vdd pdrv2 pdrv2 out out vdd out vdd vdd pdrv2 vdd pdrv2 pdrv2 pdrv2 vdd pdrv2
+ pdrv2 pdrv2 vdd pdrv2 pdrv2 out pdrv2 pdrv2 vdd out pdrv2 out out vdd out pdrv2
+ pdrv2 out vdd pdrv2 out vdd pdrv2 out out pdrv2 vdd pdrv2 out out pdrv2 out pdrv2
+ pdrv2 vdd pdrv2 out pdrv2 pdrv2 vdd pdrv2 vdd vdd vdd vdd out out out pdrv2 out
+ pdrv2 pdrv2 pdrv2 vdd pdrv2 pdrv2 pdrv2 out out pdrv2 vdd vdd out pdrv2 vdd vdd
+ vdd out out out pdrv2 pdrv2 vdd out vdd pdrv2 pdrv2 out pdrv2 out out vdd vdd pdrv2
+ pdrv2 out pdrv2 pdrv2 vdd out out pdrv2 vdd vdd out pdrv2 vdd vdd out vdd out vdd
+ pdrv2 out vdd pdrv2 pdrv2 pdrv2 vdd vdd out pdrv2 out pdrv2 out out out out pdrv2
+ vdd pdrv2 pdrv2 pdrv2 out pdrv2 out pdrv2 pdrv2 out pdrv2 vdd vdd pdrv2 vdd out
+ pdrv2 vdd vdd vdd vdd out out vdd pdrv2 out pdrv2 out pdrv2 pdrv2 pdrv2 vdd pdrv2
+ pdrv2 out pdrv2 pdrv2 pdrv2 pdrv2 vdd vdd vdd vdd out pdrv2 out vdd vdd pdrv2 pdrv2
+ out out pdrv2 vdd vdd out pdrv2 pdrv2 pdrv2 pdrv2 out pdrv2 pdrv2 out pdrv2 vdd
+ vdd out pdrv2 pdrv2 out vdd out pdrv2 vdd out out pdrv2 pdrv2 pdrv2 pdrv2 vdd pdrv2
+ pdrv2 pdrv2 out pdrv2 pdrv2 vdd pdrv2 vdd pdrv2 pdrv2 out pdrv2 out vdd pdrv2 out
+ out vdd vdd pdrv2 pdrv2 pdrv2 vdd out pdrv2 pdrv2 pdrv2 pdrv2 vdd out pdrv2 vdd
+ out out pdrv2 vdd pdrv2 out out vdd pdrv2 pdrv2 vdd pdrv2 pdrv2 pdrv2 pdrv2 out
+ pdrv2 vdd pdrv2 pdrv2 pdrv2 pdrv2 out pdrv2 pdrv2 pdrv2 vdd out pdrv2 vdd vdd out
+ out pdrv2 pdrv2 vdd vdd pdrv2 pdrv2 vdd pdrv2 pdrv2 pdrv2 pdrv2 out vdd pdrv2 out
+ pdrv2 out pdrv2 vdd out pdrv2 out pdrv2 out pdrv2 vdd out vdd pdrv2 out out pdrv2
+ pdrv2 pdrv2 pdrv2 pdrv2 pdrv2 pdrv2 vdd pdrv2 pdrv2 pdrv2 vdd pdrv2 out pdrv2 vdd
+ pdrv2 out out pdrv2 out vdd out pdrv2 pdrv2 out pdrv2 vdd pdrv2 vdd pdrv2 pdrv2
+ pdrv2 pdrv2 out pdrv2 out pdrv2 pdrv2 pdrv2 pdrv2 pdrv2 out pdrv2 vdd out pdrv2
+ pdrv2 vdd vdd out vdd pdrv2 pdrv2 vdd pdrv2 pdrv2 out pdrv2 pdrv2 pdrv2 pdrv2 vdd
+ pdrv2 pdrv2 vdd out sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT
XXM30 vss vss m1_n523_n317# m1_n523_n317# sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
XXM10 nbias vss nbias vss nbias vss vss nbias nbias nbias sky130_fd_pr__nfet_g5v0d10v5_H7BQ24
XXM22 ndrv ndrv vss ndrv vss ndrv ndrv vss vss ndrv vss ndrv out out ndrv ndrv out
+ out out vss vss ndrv vss out ndrv vss out ndrv vss ndrv ndrv ndrv ndrv out ndrv
+ ndrv out ndrv ndrv out out ndrv out ndrv out vss vss ndrv ndrv out ndrv ndrv ndrv
+ out vss vss ndrv out ndrv vss ndrv ndrv vss ndrv ndrv ndrv ndrv out ndrv ndrv out
+ ndrv ndrv ndrv ndrv ndrv vss out out ndrv vss ndrv ndrv vss ndrv ndrv out vss out
+ vss out ndrv vss ndrv vss ndrv ndrv out ndrv ndrv ndrv ndrv ndrv vss ndrv ndrv ndrv
+ ndrv out ndrv ndrv out ndrv ndrv out vss out ndrv out ndrv vss ndrv ndrv vss vss
+ vss vss ndrv out ndrv out ndrv ndrv ndrv out ndrv ndrv ndrv out ndrv ndrv ndrv vss
+ ndrv ndrv ndrv ndrv vss ndrv vss out vss vss ndrv ndrv out ndrv out vss ndrv ndrv
+ vss out out vss ndrv out ndrv ndrv ndrv vss ndrv ndrv ndrv ndrv ndrv out vss vss
+ vss vss ndrv out out ndrv out out ndrv out out ndrv out vss ndrv vss ndrv vss out
+ vss out vss out out vss ndrv ndrv ndrv out out vss out ndrv vss ndrv ndrv vss out
+ out vss out vss ndrv out ndrv ndrv ndrv vss vss ndrv vss out vss ndrv ndrv out vss
+ ndrv out out vss out vss ndrv ndrv sky130_fd_pr__nfet_g5v0d10v5_UC3VEF
.ends

.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 VGND VPWR A X VNB VPB LVPWR
X0 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=2.71875e+12p pd=2.345e+07u as=1.2375e+12p ps=1.065e+07u w=1.5e+06u l=500000u
X1 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2 X a_1711_885# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=8.13e+11p ps=7.01e+06u w=1.5e+06u l=500000u
X3 X a_1711_885# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X4 VGND A a_404_1133# VNB sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X5 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X6 VPWR a_1197_107# a_504_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.142e+11p ps=1.99e+06u w=420000u l=1e+06u
X7 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X8 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X9 a_772_151# a_404_1133# VGND VNB sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X10 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X11 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X12 LVPWR A a_404_1133# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=2.352e+11p pd=2.24e+06u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X13 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X14 VPWR a_504_1221# a_1711_885# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X15 VGND a_504_1221# a_1711_885# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X16 VGND a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X17 a_772_151# a_404_1133# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X18 a_1197_107# a_772_151# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X19 VPWR a_504_1221# a_1197_107# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=1e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCAG9S c1_n550_n500# m3_n650_n600#
X0 c1_n550_n500# m3_n650_n600# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_VCAE9S c2_n751_n500# m4_n851_n600#
X0 c2_n751_n500# m4_n851_n600# sky130_fd_pr__cap_mim_m3_2 l=5e+06u w=5e+06u
.ends

.subckt hold_cap_array holdval vss
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_1[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_2[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_3[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_4[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_5[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_6[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_6[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_6[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_6[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_6[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_6[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_6[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_6[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_7[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_7[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_7[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_7[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_7[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_7[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_7[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_7[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_8[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_8[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_8[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_8[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_8[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_8[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_8[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_8[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXC2[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
XXC2[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_9[0] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_9[1] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_9[2] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_9[3] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_9[4] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_9[5] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_9[6] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_9[7] holdval vss sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_0[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_1[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_2[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_3[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_4[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_5[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_5[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_5[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_5[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_5[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_5[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_5[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_5[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_6[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_6[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_6[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_6[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_6[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_6[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_6[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_6[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_7[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_7[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_7[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_7[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_7[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_7[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_7[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_7[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_8[0] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_8[1] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_8[2] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_8[3] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_8[4] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_8[5] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_8[6] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
Xsky130_fd_pr__cap_mim_m3_2_VCAE9S_8[7] vss holdval sky130_fd_pr__cap_mim_m3_2_VCAE9S
.ends

.subckt sample_and_hold out vdd hold in dvdd dvss ena vss
Xx1 x1/hold x3/in x1/in vdd vss balanced_switch
Xx3 vdd x3/in out ena vss follower_amp
Xx2 vdd in x1/in ena vss follower_amp
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 dvss vdd hold x1/hold dvss vdd dvdd sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_pr__diode_pw2nd_05v5_L93GHW_0 dvss hold sky130_fd_pr__diode_pw2nd_05v5_L93GHW
Xhold_cap_array_0 x3/in vss hold_cap_array
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 X A VGND VPWR VNB VPB LVPWR
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=1.113e+11p pd=1.37e+06u as=2.394e+11p ps=2.82e+06u w=420000u l=500000u
X1 VGND a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=1.7205e+12p pd=1.522e+07u as=1.197e+11p ps=1.41e+06u w=420000u l=500000u
X2 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=6.075e+11p ps=6.12e+06u w=750000u l=500000u
X3 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=6.075e+11p pd=6.12e+06u as=0p ps=0u w=750000u l=500000u
X5 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.197e+11p ps=1.41e+06u w=420000u l=500000u
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=6.104e+11p pd=5.57e+06u as=2.968e+11p ps=2.77e+06u w=1.12e+06u l=150000u
X11 VGND a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=1.961e+11p pd=2.01e+06u as=1.961e+11p ps=2.01e+06u w=740000u l=150000u
X12 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.968e+11p ps=2.77e+06u w=1.12e+06u l=150000u
X14 a_30_207# a_30_1337# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=500000u
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=2.968e+11p pd=2.77e+06u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt comparator_bias VBP VBN VDD VSS
X0 a_508011_646777# a_512471_646247# VSS sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X1 VSS VSS VBP VSS sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.232e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=2e+06u
X2 a_508011_646777# a_512471_647307# VSS sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X3 VSS VSS a_513709_648116# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=2e+06u
X4 VDD VBP VBP VDD sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.232e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=2e+06u
X5 a_508011_647837# a_512471_648367# VSS sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X6 a_508011_646247# a_512471_646247# VSS sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X7 a_508013_648897# a_512471_648367# VSS sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X8 a_513709_648116# a_508011_646247# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+12p pd=2.116e+07u as=0p ps=0u w=5e+06u l=2e+06u
X9 VBP VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X10 VBN a_513709_648116# a_508011_646247# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=3.19e+12p pd=2.374e+07u as=4.64e+12p ps=3.432e+07u w=5e+06u l=2e+06u
X11 a_513709_648116# a_508011_646247# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X12 VBN a_513709_648116# a_508011_646247# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X13 VSS VBN VBN VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=2e+06u
X14 VDD a_508011_646247# a_513709_648116# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X15 VDD a_508011_646247# a_513709_648116# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X16 a_508013_648897# VDD VSS sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X17 a_508011_646247# a_513709_648116# VBN VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X18 a_508011_646247# a_513709_648116# VBN VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X19 VBN VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X20 a_513709_648116# VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X21 a_508011_647837# a_512471_647307# VSS sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X22 VBN VBN a_508011_646247# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1.5e+07u
.ends

.subckt comparator VBP VBN VINP VINM VDD VSS VOUT
X0 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.755e+13p pd=2.0102e+08u as=0p ps=0u w=5e+06u l=2e+06u
X1 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+13p pd=2.1102e+08u as=0p ps=0u w=5e+06u l=2e+06u
X2 VSS a_512178_643337# a_512178_640243# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+12p ps=2.116e+07u w=5e+06u l=2e+06u
X3 VOUT a_515760_641405# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=2e+06u
X4 a_509030_644406# a_509030_644406# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=2e+06u
X5 VOUT a_515760_641405# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=0p ps=0u w=1e+07u l=2e+06u
X6 a_512178_640243# a_512178_643337# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X7 a_509030_644406# VINM a_508972_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+12p pd=2.116e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=2e+06u
X8 VSS a_509030_640217# a_509430_640243# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=2e+06u
X9 a_509030_640217# VINM a_508972_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+12p pd=2.116e+07u as=8.7e+12p ps=6.348e+07u w=5e+06u l=2e+06u
X10 a_512178_640243# a_509430_644503# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X11 a_512178_643337# a_512178_643337# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=2e+06u
X12 VDD a_512178_641405# a_512178_640243# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+12p ps=2.116e+07u w=5e+06u l=2e+06u
X13 a_512178_640243# a_512178_641405# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X14 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X15 VDD a_509030_644406# a_509430_644503# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=2e+06u
X16 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X17 VSS a_509430_644503# a_512178_640243# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X18 a_512178_640243# a_509430_640243# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X19 VDD VDD a_508972_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X20 VSS VSS a_508972_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X21 VSS a_512178_643337# a_512178_643337# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X22 a_512178_641405# a_512178_641405# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=2e+06u
X23 a_508972_641405# VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X24 a_508972_643337# VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X25 a_512178_641405# VINP a_508972_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+12p pd=2.116e+07u as=0p ps=0u w=5e+06u l=2e+06u
X26 a_512178_643337# VINP a_508972_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+12p pd=2.116e+07u as=0p ps=0u w=5e+06u l=2e+06u
X27 a_512178_641405# VINP a_508972_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X28 a_512178_643337# VINP a_508972_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X29 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X30 VDD a_509430_640243# a_512178_640243# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X31 a_509430_644503# a_509430_644503# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=2e+06u
X32 VDD a_512178_641405# a_512178_641405# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X33 a_508972_643337# VINP a_512178_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X34 a_508972_641405# VINP a_512178_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X35 a_508972_641405# VINP a_512178_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X36 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X37 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X38 a_508972_643337# VINP a_512178_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X39 a_509430_640243# a_509030_640217# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X40 VSS a_509030_640217# a_509030_640217# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=2e+06u
X41 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X42 VSS a_509430_644503# a_509430_644503# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X43 a_509430_640243# a_509430_640243# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=2e+06u
X44 a_508972_641405# VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X45 a_508972_643337# VBP VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X46 a_509030_640217# VINM a_508972_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X47 a_509030_644406# VINM a_508972_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X48 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X49 VSS a_512178_640243# a_515760_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=2e+06u
X50 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X51 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X52 VDD a_512178_640243# a_515760_641405# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u l=2e+06u
X53 a_509430_644503# a_509030_644406# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X54 VDD a_509030_644406# a_509030_644406# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X55 VDD a_509430_640243# a_509430_640243# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X56 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X57 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X58 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X59 VSS VBN a_508972_641405# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X60 a_508972_641405# VINM a_509030_644406# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X61 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X62 a_509030_640217# a_509030_640217# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X63 VDD VBP a_508972_643337# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X64 a_508972_643337# VINM a_509030_640217# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X65 a_508972_641405# VINM a_509030_644406# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X66 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X67 a_508972_643337# VINM a_509030_640217# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
.ends

.subckt comparator_top VINM VINP VDD VOUT DVDD DVSS VSS
Xsky130_fd_sc_hvl__lsbufhv2lv_1_0 VOUT comparator_0/VOUT DVSS VDD DVSS VDD DVDD sky130_fd_sc_hvl__lsbufhv2lv_1
Xcomparator_bias_0 comparator_0/VBP comparator_0/VBN VDD VSS comparator_bias
Xcomparator_0 comparator_0/VBP comparator_0/VBN VINP VINM VDD VSS comparator_0/VOUT
+ comparator
.ends

.subckt EF_ADCS0808NSCM hold ena cmp dac_out vhigh vlow b0 b1 b2 b3 b4 b5 b6 b7 inp[0]
+ inp[1] inp[2] inp[3] inp[4] inp[5] inp[6] inp[7] in[0] in[1] in[2] dvdd vss vdd
+ dvss
Xsample_and_hold_0 sample_and_hold_0/out vdd hold sbamuxm4_0/muxout dvdd dvss ena
+ vss sample_and_hold
Xcomparator_top_0 dac_out sample_and_hold_0/out vdd cmp dvdd dvss vss comparator_top
X0 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=1.49466e+14p pd=1.30757e+09u as=1.624e+13p ps=1.352e+08u w=1e+06u l=1e+06u
X1 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=1.66026e+14p pd=1.49016e+09u as=0p ps=0u w=1e+06u l=1e+06u
X2 dac_3v_column_0[0].out1_0_1 dac_3v_8bit_0/b0a a_25577_n4028# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=6.09e+13p pd=5.418e+08u as=2.65986e+14p ps=2.29124e+09u w=1e+06u l=500000u
X4 a_25384_n7619# dac_3v_8bit_0/b0b dac_3v_column_0[2].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X5 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
D0 dvss b5 sky130_fd_pr__diode_pw2nd_05v5
X6 a_21663_n2566# vss a_21663_n2566# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X7 a_26184_n2566# vss a_25577_n2963# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X8 a_31412_n17214# dac_3v_8bit_0/b0a dac_3v_column_odd_0[6].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X9 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbp dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=2.064e+07u as=0p ps=0u w=1e+06u l=1e+06u
X10 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n55353_n19355# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X11 a_n27017_n925# a_n25859_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X12 dac_3v_column_odd_0[0].out1_0_3 dac_3v_8bit_0/b0a a_31605_n5095# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X13 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X14 dac_3v_8bit_0/b1b dac_3v_8bit_0/b1a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X15 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X a_n53983_n17697# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X16 a_20024_n2963# a_20863_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X17 a_21663_n20686# vss a_20863_n20410# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X18 dac_3v_column_odd_0[2].out1_0_0 dac_3v_8bit_0/b0b a_22563_n9359# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X19 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X20 a_24070_n17887# a_25577_n17887# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X21 a_29905_n18279# a_31412_n18279# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X22 dac_3v_column_odd_0[4].res_in0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[4].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X23 a_n54937_n18785# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n54657_n18785# dvdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X24 dvss bias_0.bi__pmirr_0.gate_cas dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X25 dvdd a_n53523_n22049# testbuffer_0.tb__mux_0.tbm__passgate_5.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X26 dac_3v_column_0[7].out1_0_3 dac_3v_8bit_0/b0a a_30098_n18952# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X27 a_31412_n16147# dac_3v_column_odd_0[5].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X28 a_33719_n14291# vdd dac_3v_column_odd_0[5].res_in0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X29 dvss level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b3a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=5.29492e+13p pd=4.7763e+08u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X30 dac_3v_8bit_0/b4b dac_3v_8bit_0/b4a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X31 dvss dac_3v_8bit_0/b3a dac_3v_8bit_0/b3b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X32 dac_3v_column_odd_0[0].out1_0_0 dac_3v_8bit_0/b0a a_22563_n5095# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X33 a_28398_n2290# a_29905_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X34 dac_3v_column_odd_0[3].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_odd_0[3].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X35 a_20156_n11094# vdd dac_3v_column_odd_0[3].dum_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X36 testbuffer_0.tb__mux_0.tbm__passgate_3.en a_n54301_n18241# dvss dvss sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X37 a_30098_n9359# a_31605_n9359# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X38 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=7.31448e+13p pd=6.16795e+08u as=1.827e+13p ps=1.6254e+08u w=1e+06u l=500000u
X39 dac_3v_column_odd_0[3].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[3].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X40 a_20156_n10027# vss a_20156_n10027# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X41 sbamuxm4_0/vb[5] a_n32029_7560# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X42 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X43 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=4.06e+12p pd=3.612e+07u as=6.38e+12p ps=5.676e+07u w=1e+06u l=4e+06u
X44 a_30705_n20686# vss a_30705_n20686# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X45 a_29905_n7619# dac_3v_8bit_0/b0a dac_3v_column_0[2].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X46 dac_3v_column_odd_0[4].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_odd_0[4].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X47 dac_3v_column_odd_0[3].dum_in0 vss a_34426_n11252# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X48 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X49 a_20156_n19622# vdd a_20156_n19622# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X50 a_28398_n19346# dac_3v_8bit_0/b0a dac_3v_column_odd_0[7].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X51 a_23170_n12950# dac_3v_8bit_0/b2a dac_3v_column_odd_0[4].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X52 dac_3v_column_odd_0[1].out1_0_2 dac_3v_8bit_0/b0b a_28591_n7227# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X53 dac_3v_8bit_0/b0a dac_3v_8bit_0/b0b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X54 a_23877_n19346# dac_3v_8bit_0/b0a dac_3v_column_odd_0[7].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X55 a_28686_3107# b3 dvss dvss sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X56 dac_3v_column_0[1].dum1_in dac_3v_column_0[1].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X57 a_20863_n8053# vss a_20863_n8053# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X58 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X59 sbamuxm4_0/ibn[1] bias_0.bi__pmirr_0.gate_cas a_n41084_7586# dvss sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=2.064e+07u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X60 dac_3v_column_0[6].out_3 dac_3v_8bit_0/b3b dac_3v_column_0[6].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X61 a_28591_n10424# a_30098_n10424# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X62 dvss a_27058_3107# a_27058_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.2375e+12p ps=1.065e+07u w=1.5e+06u l=500000u
X63 dac_3v_8bit_0/b0b level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=8.4e+11p pd=8.24e+06u as=0p ps=0u w=750000u l=500000u
X64 dac_3v_column_0[6].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_0[6].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X65 a_20156_n15358# vss dac_3v_column_odd_0[5].dum_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X66 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X67 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X68 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=4.06e+12p pd=3.612e+07u as=6.38e+12p ps=5.676e+07u w=1e+06u l=4e+06u
X69 dvss dac_3v_8bit_0/b4a dac_3v_8bit_0/b4b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X70 vdd level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b2a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.68e+12p ps=1.424e+07u w=1.5e+06u l=500000u
X71 a_31412_n2290# a_32919_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X72 dac_3v_column_0[1].out1_0_0 dac_3v_8bit_0/b0b a_22563_n6160# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X73 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X74 a_29905_n14015# dac_3v_8bit_0/b0a dac_3v_column_0[5].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X75 dac_3v_column_0[5].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[5].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X76 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X77 a_22370_n18279# dac_3v_8bit_0/b0a dac_3v_column_0[7].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X78 a_n55646_9265# a_n55646_9265# dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X79 dvss a_28686_3107# a_28686_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.2375e+12p ps=1.065e+07u w=1.5e+06u l=500000u
X80 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X81 a_22752_2837# a_23114_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X82 a_n53523_n22049# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._17_.X dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X83 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X84 dvdd a_22174_3107# a_23114_3404# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X85 a_22370_n2290# a_23877_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X86 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X87 dvss level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b4a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X88 dac_3v_column_0[4].out1_0_1 dac_3v_8bit_0/b0a a_25577_n12556# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X89 a_20156_n7895# vdd dac_3v_column_0[2].dum1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X90 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X91 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X92 testbuffer_0.tb__mux_0.tbm__passgate_0.en a_n54221_n16635# dvss dvss sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X93 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X94 a_22370_n11883# a_23877_n11883# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X95 dvss bias_0.bi__nmirr_0.gate_n a_n42000_9346# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X96 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbn dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.61e+12p pd=2.322e+07u as=0p ps=0u w=1e+06u l=500000u
X97 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X98 dvss level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4.2e+11p ps=4.12e+06u w=750000u l=500000u
X99 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X100 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n53615_n20961# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u
X101 a_34426_n16581# vss a_34426_n16581# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X102 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X103 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=1.856e+13p pd=1.4076e+08u as=0p ps=0u w=1e+06u l=1e+06u
X104 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n48623_n15278# inp[1] dvdd sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=2.064e+07u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X105 dac_3v_column_0[6].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[6].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X106 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=8.12e+12p pd=6.412e+07u as=0p ps=0u w=2e+06u l=4e+06u
X107 a_33719_n3631# vss a_33719_n3631# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X108 dac_3v_column_odd_0[2].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[2].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X109 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X110 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X111 a_23877_n3355# a_25384_n3355# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X112 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X113 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.432e+07u as=0p ps=0u w=4e+06u l=1e+06u
X114 dac_3v_8bit_0/b2b dac_3v_8bit_0/b2a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=8.4e+11p pd=8.24e+06u as=0p ps=0u w=750000u l=500000u
X115 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X116 a_25384_n6554# a_26891_n6554# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X117 a_30098_n12556# a_31605_n12556# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X118 dac_3v_column_0[3].dum1_in dac_3v_column_0[3].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X119 dvss bias_0.bi__nmirr_0.gate_n dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X120 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n47185_n21248# inp[4] dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X121 dac_3v_column_odd_0[4].out1_0_0 dac_3v_8bit_0/b0a a_22563_n13623# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X122 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X123 dac_3v_column_odd_0[4].out_3 dac_3v_8bit_0/b3a dac_3v_column_odd_0[4].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X124 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.64e+12p ps=4.128e+07u w=1e+06u l=1e+06u
X125 dac_3v_column_odd_0[3].in_5 vss dac_3v_column_odd_0[3].in_5 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=500000u
X126 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X127 dvdd bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbp dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.32e+12p ps=2.064e+07u w=1e+06u l=1e+06u
X128 vdd dac_3v_8bit_0/b2a dac_3v_8bit_0/b2b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.68e+12p ps=1.424e+07u w=1.5e+06u l=500000u
X129 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=1.624e+13p pd=1.352e+08u as=0p ps=0u w=1e+06u l=1e+06u
X130 dac_3v_column_odd_0[0].dum_in0 vss a_34426_n4856# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X131 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X132 sbamuxm4_0/vb[3] a_n32029_10092# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X133 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X134 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X135 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X136 a_33719_n14291# vss dac_3v_column_odd_0[5].res_in0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X137 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X138 dvss level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.1e+11p ps=2.06e+06u w=750000u l=500000u
X139 sbamuxm4_0/ibp[3] bias_0.bi__pmirr_0.gate a_n42353_12567# dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=3.16e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X140 a_n55233_n20443# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output8.A dvss dvss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X141 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X142 a_n55858_5903# a_n55858_8035# dvss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X143 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X144 vdd dac_3v_8bit_0/b7b dac_3v_8bit_0/b7a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.68e+12p ps=1.424e+07u w=1.5e+06u l=500000u
X145 dac_3v_8bit_0/b6b level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X146 a_26891_n9751# dac_3v_8bit_0/b0b dac_3v_column_0[3].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X147 a_n54427_5925# dvss dvss sky130_fd_pr__res_xhigh_po w=350000u l=7e+06u
X148 dvss level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4.2e+11p ps=4.12e+06u w=750000u l=500000u
X149 a_26891_n5487# dac_3v_8bit_0/b0a dac_3v_column_0[1].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X150 a_25577_n18952# a_27084_n18952# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X151 dvss a_24742_3404# a_24380_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.2375e+12p ps=1.065e+07u w=1.5e+06u l=500000u
X152 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X153 dac_3v_column_odd_0[4].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_odd_0[4].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X154 a_25384_n4422# dac_3v_8bit_0/b0b dac_3v_column_odd_0[0].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X155 dvss a_n54035_n19757# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output5.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X156 follower_amp_0.vcomn1 dac_out a_14987_n11444# vss sky130_fd_pr__nfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X157 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X158 dac_3v_column_0[4].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_0[4].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X159 dac_3v_column_0[3].out0_2 dac_3v_8bit_0/b3a dac_3v_column_0[3].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X160 a_n26631_n925# a_n27789_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X161 bias_0.bi__amplifier_0.inn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvdd dvdd sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=1e+06u
X162 dac_3v_column_0[0].out1_0_3 dac_3v_8bit_0/b0b a_31605_n4028# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X163 a_20863_n12317# vss a_20863_n12317# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X164 dac_3v_column_0[0].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[0].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X165 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.832e+07u as=9.28e+12p ps=7.328e+07u w=2e+06u l=4e+06u
X166 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X167 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X168 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X169 dac_3v_column_odd_0[1].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_odd_0[1].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X170 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X171 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X172 dac_3v_column_odd_0[3].out1_0_0 dac_3v_8bit_0/b0b a_22563_n11491# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X173 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X174 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X175 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X a_n55547_n16609# dvss dvss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X176 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._19_.X a_n53289_n21505# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X177 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X178 dac_3v_column_odd_0[7].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_odd_0[7].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X179 dac_3v_column_0[5].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[5].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X180 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X181 a_31412_n12950# dac_3v_column_odd_0[4].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X182 dac_3v_column_odd_0[1].res_in1 vdd a_20863_n6988# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X183 a_20863_n2290# vss a_20863_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X184 dvss level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b5a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X185 a_23170_n19346# dac_3v_8bit_0/b1a dac_3v_column_odd_0[7].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X186 a_32919_n2724# vdd a_32919_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X187 sbamuxm4_0/vb[6] a_n32029_6716# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X188 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X189 level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=4.2e+11p pd=4.12e+06u as=0p ps=0u w=750000u l=500000u
X190 dac_3v_column_0[1].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[1].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X191 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X192 dac_3v_8bit_0/out_unbuf dac_3v_8bit_0/b7b dac_3v_column_odd_0[2].in_5 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X193 a_29905_n4422# dac_3v_8bit_0/b0a dac_3v_column_odd_0[0].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X194 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.64e+12p ps=4.128e+07u w=1e+06u l=1e+06u
X195 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X196 dac_3v_column_0[6].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_0[6].res1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X197 a_n54691_n21255# a_n54441_n21531# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output8.A dvdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X198 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X199 a_33719_n2566# vdd vhigh vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X200 a_n32750_1515# a_n31275_1643# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X201 dac_3v_column_0[2].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_0[2].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X202 dac_3v_8bit_0/b3b dac_3v_8bit_0/b3a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X203 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X204 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X205 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X206 a_23877_n2724# vdd a_23877_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X207 dac_3v_column_odd_0[4].out4 dac_3v_8bit_0/b4b dac_3v_column_0[4].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X208 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X209 a_n42000_7938# bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[0] dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.32e+12p ps=2.064e+07u w=1e+06u l=2e+06u
X210 a_n40589_11671# bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.gate_cas dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=3.16e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X211 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X212 dac_3v_column_0[6].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[6].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X213 a_22370_n7619# dac_3v_8bit_0/b0a dac_3v_column_0[2].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X214 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X215 a_28398_n15082# a_29905_n15082# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X216 dvss a_25430_3107# a_25430_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.2375e+12p ps=1.065e+07u w=1.5e+06u l=500000u
X217 a_20156_n2566# vdd a_20156_n2566# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X218 a_24677_n2566# vdd a_24070_n2963# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X219 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X220 vdd dac_3v_8bit_0/b0b dac_3v_8bit_0/b0a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X221 vdd a_23802_2206# level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X222 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C a_n53615_n20961# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X223 vdd level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=7.12e+06u w=1.5e+06u l=500000u
X224 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X225 a_30314_2371# a_30314_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X226 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X227 a_22370_n15082# dac_3v_8bit_0/b0a dac_3v_column_odd_0[5].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X228 dvss in[0] a_n55547_n16609# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X229 follower_amp_0.nbias follower_amp_0.nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X230 dac_3v_column_0[7].out1_0_1 dac_3v_8bit_0/b0b a_24070_n18952# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X231 dac_3v_column_0[4].out1_0_2 dac_3v_8bit_0/b0b a_28591_n12556# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X232 bias_0.bi__amplifier_0.diff bias_0.bi__amplifier_0.inn bias_0.bi__pmirr_0.gate dvss sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=1.264e+07u as=5.8e+11p ps=6.32e+06u w=500000u l=8e+06u
X233 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X234 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X235 a_28686_2206# a_28686_2371# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X236 a_30098_n2963# a_31605_n2963# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X237 dac_3v_column_odd_0[6].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_odd_0[6].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X238 a_28398_n20844# vss a_28398_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X239 a_26891_n18279# dac_3v_8bit_0/b0b dac_3v_column_0[7].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X240 dvss a_n54345_n20265# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.X dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X241 a_34426_n13384# vdd a_34426_n13384# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X242 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=9.28e+12p pd=8.256e+07u as=9.28e+12p ps=8.256e+07u w=1e+06u l=500000u
X243 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X244 a_22370_n18279# dac_3v_8bit_0/b0b dac_3v_column_0[7].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X245 dac_3v_column_odd_0[7].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[7].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X246 a_24677_n20686# vdd a_24677_n20686# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X247 dac_3v_column_0[2].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_0[2].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X248 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X249 dvss level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b7b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X250 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X251 a_31412_n14015# dac_3v_8bit_0/b0a dac_3v_column_0[5].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X252 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X253 level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X254 a_27691_n2566# vss a_27084_n2963# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X255 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X256 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X257 a_23170_n17214# dac_3v_8bit_0/b1a dac_3v_column_odd_0[6].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
D1 dvss b4 sky130_fd_pr__diode_pw2nd_05v5
X258 level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=4.2e+11p pd=4.12e+06u as=0p ps=0u w=750000u l=500000u
X259 a_24070_n14688# a_25577_n14688# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X260 dac_3v_column_odd_0[6].out1_0_2 dac_3v_8bit_0/b0b a_27084_n17887# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X261 dac_3v_column_odd_0[2].out1_0_1 dac_3v_8bit_0/b0a a_24070_n9359# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X262 dac_3v_column_0[2].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[2].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X263 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.58e+07u as=1.74e+12p ps=1.548e+07u w=1e+06u l=4e+06u
X264 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X265 dvss bias_0.bi__pmirr_0.gate_cas dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X266 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X267 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X268 dac_3v_column_odd_0[7].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[7].res_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X269 dac_3v_column_odd_0[4].out1_0_1 dac_3v_8bit_0/b0b a_25577_n13623# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X270 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X271 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X272 a_30098_n20019# a_31605_n20019# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X273 bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__pmirr_0.vbn dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X274 a_26891_n4422# a_28398_n4422# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X275 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X276 a_30098_n6160# a_31605_n6160# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X277 dac_3v_column_0[2].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_0[2].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X278 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X279 a_22370_n11883# dac_3v_8bit_0/b0a dac_3v_column_0[4].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X280 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X281 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X282 dac_3v_column_odd_0[2].out_5 dac_3v_8bit_0/b5a dac_3v_column_odd_0[3].out4 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X283 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n46909_n21248# inp[4] dvss sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=2.064e+07u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X284 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X285 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X286 a_28398_n16147# dac_3v_8bit_0/b0a dac_3v_column_0[6].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X287 a_20156_n16423# vdd a_20156_n16423# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X288 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X289 dvss a_n54443_n22593# testbuffer_0.tb__mux_0.tbm__passgate_6.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X290 a_29905_n17214# a_31412_n17214# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X291 dac_3v_column_odd_0[5].dum_in1 dac_3v_column_odd_0[5].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X292 dac_3v_column_odd_0[6].dum_out1 vss a_34426_n18713# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X293 a_23877_n16147# dac_3v_8bit_0/b0a dac_3v_column_0[6].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X294 a_n42000_7586# bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[1] dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X295 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X296 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.432e+07u as=0p ps=0u w=4e+06u l=1e+06u
X297 a_26008_2837# a_25430_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=1e+06u
X298 dac_3v_column_odd_0[1].out1_0_3 dac_3v_8bit_0/b0b a_30098_n7227# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X299 a_25384_n19346# a_26891_n19346# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X300 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X301 dac_3v_column_odd_0[5].res_in1 a_22563_n15755# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X302 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X303 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n48347_n18263# inp[2] dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X304 a_31605_n17887# dac_3v_column_odd_0[6].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X305 a_23802_2371# a_24380_2837# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.142e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=1e+06u
X306 dac_3v_column_0[2].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_0[2].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X307 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X308 vdd level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b1a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.68e+12p ps=1.424e+07u w=1.5e+06u l=500000u
X309 a_20156_n12159# vss dac_3v_column_0[4].dum1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X310 a_20863_n6988# vdd a_20863_n6988# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X311 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X312 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X313 a_23877_n20844# vdd a_23877_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X314 a_20863_n17648# vdd a_20863_n17648# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X315 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X316 a_29905_n8686# dac_3v_8bit_0/b0b dac_3v_column_odd_0[2].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X317 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=1.45e+12p pd=1.29e+07u as=0p ps=0u w=1e+06u l=4e+06u
X318 a_27636_2837# a_27998_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X319 dac_3v_column_0[1].out1_0_1 dac_3v_8bit_0/b0a a_24070_n6160# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X320 a_33719_n19622# vdd vlow vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X321 dac_3v_column_odd_0[1].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[1].res_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X322 dvdd bias_basis_current_0.bb__pmirr_0.vbp bias_0.bi__amplifier_0.bias dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=1e+06u
X323 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X324 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X325 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n46909_n24233# inp[7] dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X326 dac_3v_column_odd_0[3].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_odd_0[3].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X327 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X328 dvss a_n55547_n19873# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X329 a_30314_3107# b2 dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X330 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X331 dac_3v_8bit_0/b7a dac_3v_8bit_0/b7b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X332 a_25384_n17214# dac_3v_8bit_0/b0a dac_3v_column_odd_0[6].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X333 dac_3v_column_odd_0[6].res_in1 vss a_20863_n17648# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X334 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X335 a_24380_2837# a_24742_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X336 dvss a_27998_3404# a_27636_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X337 vdd level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=7.12e+06u w=1.5e+06u l=500000u
X338 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X339 a_31412_n19346# dac_3v_8bit_0/b0b dac_3v_column_odd_0[7].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X340 a_21663_n20686# vdd a_20863_n20410# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X341 dvdd a_23802_3107# a_24742_3404# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X342 dvss a_n53983_n17697# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X343 a_23877_n7619# a_25384_n7619# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X344 dvdd a_n54443_n22593# testbuffer_0.tb__mux_0.tbm__passgate_6.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X345 dvss dac_3v_8bit_0/b1a dac_3v_8bit_0/b1b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X346 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X347 dac_3v_column_odd_0[3].out1_0_2 dac_3v_8bit_0/b0a a_27084_n11491# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X348 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X349 a_n54443_n22593# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.X dvss dvss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X350 a_25384_n16147# a_26891_n16147# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X351 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X352 dac_3v_column_odd_0[2].dum_in0 vdd a_34426_n9120# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X353 dvss dac_3v_8bit_0/b4a dac_3v_8bit_0/b4b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X354 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X355 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C a_n54487_n21933# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5725e+11p ps=2.99e+06u w=420000u l=150000u
X356 dac_3v_column_0[1].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[1].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X357 dac_3v_column_odd_0[6].out4 dac_3v_8bit_0/b4b dac_3v_column_odd_0[6].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X358 dac_3v_column_odd_0[7].out0_2 dac_3v_8bit_0/b3b dac_3v_column_odd_0[7].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X359 dac_3v_column_odd_0[5].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[5].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X360 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvss sky130_fd_pr__nfet_01v8_lvt ad=1.044e+13p pd=8.476e+07u as=2.32e+12p ps=1.832e+07u w=2e+06u l=1e+06u
X361 a_27084_n16820# a_28591_n16820# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X362 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X363 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbp dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X364 dac_3v_column_odd_0[0].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_odd_0[0].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X365 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X366 dac_3v_column_odd_0[7].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[7].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X367 a_28398_n10818# dac_3v_8bit_0/b0b dac_3v_column_odd_0[3].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X368 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X369 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X370 a_23170_n12950# dac_3v_8bit_0/b2b dac_3v_column_odd_0[4].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X371 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._07_.X a_n55313_n22049# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X372 bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas dvss sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=2.064e+07u as=0p ps=0u w=1e+06u l=2e+06u
X373 dac_3v_column_0[0].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[0].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X374 a_25384_n8686# dac_3v_8bit_0/b0a dac_3v_column_odd_0[2].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X375 a_25384_n3355# a_26891_n3355# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X376 a_22370_n4422# dac_3v_8bit_0/b0a dac_3v_column_odd_0[0].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X377 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X378 dac_3v_8bit_0/b6b level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=8.4e+11p pd=8.24e+06u as=0p ps=0u w=750000u l=500000u
X379 vdd level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b3a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.68e+12p ps=1.424e+07u w=1.5e+06u l=500000u
X380 dac_3v_column_0[3].out1_0_0 dac_3v_8bit_0/b0a a_22563_n10424# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X381 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X382 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X383 a_28398_n2290# vss a_28398_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X384 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X385 dac_3v_column_odd_0[6].res_in0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[6].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X386 dac_3v_column_odd_0[6].res_in0 dac_3v_column_odd_0[6].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X387 dac_3v_column_0[3].out_3 dac_3v_8bit_0/b3a dac_3v_column_0[3].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X388 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X389 dac_3v_column_odd_0[6].out1_0_3 dac_3v_8bit_0/b0b a_30098_n17887# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X390 a_33719_n20686# vdd a_33112_n21083# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X391 a_n55547_n19873# in[1] dvss dvss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X392 dac_3v_column_odd_0[6].out1_0_1 dac_3v_8bit_0/b0a a_24070_n17887# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X393 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X394 dvss a_32882_3404# a_32520_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.2375e+12p ps=1.065e+07u w=1.5e+06u l=500000u
X395 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output5.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X396 vdd dac_3v_8bit_0/b1a dac_3v_8bit_0/b1b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X397 dac_3v_column_odd_0[6].out_5 dac_3v_8bit_0/b5a dac_3v_column_odd_0[7].out4 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X398 dac_3v_column_odd_0[4].out1_0_3 dac_3v_8bit_0/b0b a_31605_n13623# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X399 dac_3v_column_odd_0[1].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[1].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X400 dvss dvss bandgap_0.bg__pnp_group_0.eg sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=1
X401 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X402 dac_3v_8bit_0/b0b level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X403 a_n23132_n3629# a_n21227_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X404 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n53983_n17697# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X405 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X406 a_n54443_n22593# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.X dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X407 a_24070_n5095# a_25577_n5095# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X408 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X409 a_25430_2371# a_25430_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X410 a_26891_n15082# dac_3v_8bit_0/b0b dac_3v_column_odd_0[5].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X411 dvdd testbuffer_0.tb__mux_0.tbm__passgate_2.en a_n47185_n18263# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X412 dvss level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.1e+11p ps=2.06e+06u w=750000u l=500000u
X413 dac_3v_column_odd_0[0].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_odd_0[0].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X414 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X415 dac_3v_column_odd_0[6].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[6].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X416 a_n32750_455# a_n31275_n477# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X417 a_22370_n15082# dac_3v_8bit_0/b0b dac_3v_column_odd_0[5].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X418 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X419 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X a_n55527_n18241# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X420 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X421 a_34426_n3789# vdd a_34426_n3789# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X422 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X423 dac_3v_column_0[7].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[7].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X424 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X425 testbuffer_0.tb__mux_0.tbm__passgate_0.en a_n54221_n16635# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X426 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X427 a_31412_n2290# vss a_31412_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X428 dac_3v_8bit_0/b3b dac_3v_8bit_0/b3a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
D2 dvss b6 sky130_fd_pr__diode_pw2nd_05v5
X429 dac_3v_column_0[0].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_0[0].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X430 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X431 a_24070_n11491# a_25577_n11491# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X432 dac_3v_column_odd_0[2].res_out1 dac_3v_column_odd_0[2].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X433 dvss a_n55681_n22593# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X434 a_23170_n4422# dac_3v_8bit_0/b1b dac_3v_column_odd_0[0].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X435 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X436 testbuffer_0.tb__mux_0.tbm__passgate_5.en a_n53523_n22049# dvss dvss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X437 dac_3v_column_odd_0[2].out4 dac_3v_8bit_0/b4a dac_3v_column_odd_0[2].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X438 a_29905_n20410# vss a_29905_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X439 dac_3v_column_odd_0[1].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[1].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X440 sbamuxm4_0/vb[0] a_n32029_11780# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X441 level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.4e+11p pd=7.12e+06u as=0p ps=0u w=1.5e+06u l=500000u
X442 a_29905_n20844# vdd a_29905_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X443 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X444 dac_3v_column_0[6].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_0[6].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X445 dac_3v_column_0[0].res1_in vdd a_20863_n3789# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X446 dac_3v_column_0[0].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_0[0].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X447 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X448 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X449 dvdd a_n55353_n19355# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X450 follower_amp_0.vcomn2 dac_3v_8bit_0/out_unbuf follower_amp_0.pdrv2 vss sky130_fd_pr__nfet_03v3_nvt ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X451 dac_3v_column_0[6].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[6].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X452 a_23877_n10818# dac_3v_8bit_0/b0b dac_3v_column_odd_0[3].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X453 a_22370_n2290# vss a_22370_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X454 a_26891_n2724# vss a_26891_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X455 dac_3v_column_odd_0[0].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_odd_0[0].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X456 dac_3v_column_0[7].res1_in a_22370_n18279# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X457 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X458 a_33719_n19622# vss vlow vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X459 bias_0.bi__amplifier_0.mirr bias_0.bi__pmirr_0.fb bias_0.bi__amplifier_0.diff dvss sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=6.32e+06u as=0p ps=0u w=500000u l=8e+06u
X460 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X461 dac_3v_column_odd_0[0].out_5 dac_3v_8bit_0/b5a dac_3v_column_odd_0[0].out4 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X462 follower_amp_0.ndrv dac_3v_8bit_0/out_unbuf follower_amp_0.vcomp vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=1.16e+12p ps=1.032e+07u w=1e+06u l=500000u
X463 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X464 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X465 dac_3v_column_odd_0[2].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[2].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X466 a_23170_n6554# dac_3v_8bit_0/b1b dac_3v_column_odd_0[1].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X467 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output7.A a_n53197_n19329# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X468 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output5.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X469 dac_3v_column_odd_0[1].res_out1 dac_3v_8bit_0/b0b dac_3v_column_0[2].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X470 bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X471 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X472 a_22563_n21083# a_24070_n21083# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X473 a_33719_n7895# vss dac_3v_column_odd_0[2].res_in0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X474 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=1.032e+07u w=1e+06u l=4e+06u
X475 dac_3v_column_odd_0[5].dum_in0 vss a_34426_n15516# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X476 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X477 a_26891_n11883# dac_3v_8bit_0/b0b dac_3v_column_0[4].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X478 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.A a_n55681_n18241# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X479 dvss a_31942_3107# a_31942_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.2375e+12p ps=1.065e+07u w=1.5e+06u l=500000u
X480 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X481 a_22370_n11883# dac_3v_8bit_0/b0b dac_3v_column_0[4].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X482 dac_3v_column_odd_0[3].in_5 vdd dac_3v_column_odd_0[3].in_5 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X483 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X484 a_33719_n7895# vdd a_33719_n7895# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X485 bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=6.96e+12p pd=5.496e+07u as=1.74e+12p ps=1.432e+07u w=2e+06u l=4e+06u
X486 vdd level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b1a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X487 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X488 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X489 a_26891_n20410# a_28398_n20410# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X490 dvss a_30314_3107# a_30314_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X491 vdd dac_3v_8bit_0/b2a dac_3v_8bit_0/b2b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X492 a_28398_n11883# a_29905_n11883# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X493 dac_3v_column_0[3].res1_in vss a_20863_n10185# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X494 a_n40589_12119# bias_0.bi__pmirr_0.gate sbamuxm4_0/ibp[0] dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=3.16e+06u as=5.8e+11p ps=6.32e+06u w=500000u l=2e+06u
X495 dvdd a_n55681_n22593# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X496 a_23877_n7619# dac_3v_8bit_0/b0b dac_3v_column_0[2].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X497 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X498 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X499 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 dvdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.29e+07u as=5.8e+11p ps=5.16e+06u w=1e+06u l=4e+06u
X500 dac_3v_8bit_0/b0b level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X501 a_26184_n2566# vdd a_25577_n2963# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X502 a_20156_n17490# vss a_20156_n17490# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X503 dac_3v_8bit_0/b4a level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X504 dac_3v_column_odd_0[1].out4 dac_3v_8bit_0/b4b dac_3v_column_0[1].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X505 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._17_.X a_n53523_n22049# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X506 a_27058_2206# a_27058_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X507 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X508 dac_3v_column_odd_0[1].res_out1 dac_3v_column_odd_0[1].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X509 vdd a_25430_2206# level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X510 vdd level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=7.12e+06u w=1.5e+06u l=500000u
X511 dac_3v_column_0[2].out0_1_1 dac_3v_8bit_0/b2b dac_3v_column_0[2].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X512 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X513 a_n54345_n20265# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.5725e+11p pd=2.99e+06u as=0p ps=0u w=420000u l=150000u
X514 follower_amp_0.pbias follower_amp_0.nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X515 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X516 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n55353_n19355# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X517 vlow dac_3v_column_odd_0[7].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X518 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X519 dvdd a_n53615_n20961# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X520 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X521 dvss level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4.2e+11p ps=4.12e+06u w=750000u l=500000u
X522 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X523 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X524 a_n48347_n18263# a_n48623_n18263# dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X525 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X526 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X527 a_34426_n10185# vdd a_34426_n10185# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X528 dac_3v_column_odd_0[2].res_in1 a_22563_n9359# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X529 dac_3v_column_0[1].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[1].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X530 dac_3v_column_0[6].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[6].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X531 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X532 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X a_n55547_n16609# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u
X533 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X534 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X535 a_33719_n20686# vss a_33112_n21083# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X536 a_n47950_6120# bias_0.bi__amplifier_0.bias bias_0.bi__amplifier_0.diff dvss sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=6.32e+06u as=0p ps=0u w=500000u l=4e+06u
X537 dac_3v_column_odd_0[6].out1_0_3 dac_3v_8bit_0/b0a a_30098_n17887# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X538 dac_3v_column_odd_0[4].out1_0_2 dac_3v_8bit_0/b0a a_28591_n13623# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X539 dac_3v_column_odd_0[3].dum_out1 vss a_34426_n12317# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X540 a_33719_n11094# vdd a_33719_n11094# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X541 dac_3v_column_0[5].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[5].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X542 a_20156_n10027# vdd a_20156_n10027# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X543 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=9.28e+12p ps=7.328e+07u w=2e+06u l=4e+06u
X544 a_n53825_n18785# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output4.A dvdd sky130_fd_pr__pfet_01v8_hvt ad=7.9e+11p pd=7.58e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X545 a_25384_n12950# a_26891_n12950# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X546 a_20156_n8962# vss a_20156_n8962# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X547 dac_3v_column_0[2].out1_0_2 dac_3v_8bit_0/b0b a_28591_n8292# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X548 level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X549 dvss dvss bandgap_0.bg__pnp_group_0.eg sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=1
X550 dac_3v_column_0[2].out0_2 dac_3v_8bit_0/b3b dac_3v_column_0[2].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X551 dac_3v_column_odd_0[1].out1_0_2 dac_3v_8bit_0/b0a a_28591_n7227# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X552 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X553 a_27084_n13623# a_28591_n13623# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X554 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X555 dac_3v_column_0[6].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_0[6].res1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X556 dac_3v_column_0[3].out1_0_1 dac_3v_8bit_0/b0b a_25577_n10424# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X557 dac_3v_column_0[7].out1_0_3 dac_3v_8bit_0/b0a a_31605_n18952# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X558 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X559 dac_3v_column_odd_0[5].out_3 dac_3v_8bit_0/b3b dac_3v_column_odd_0[5].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X560 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X561 a_n53645_n19873# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n53925_n19873# dvdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X562 dac_3v_column_odd_0[5].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[5].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X563 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X564 dac_3v_8bit_0/b6a dac_3v_8bit_0/b6b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X565 dvss level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b2a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X566 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X567 dvss level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b5a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X568 a_32212_n20686# vdd a_32212_n20686# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X569 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X570 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n53983_n17697# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u
X571 dac_3v_column_odd_0[0].out1_0_0 dac_3v_8bit_0/b0b a_22563_n5095# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X572 dac_3v_column_odd_0[4].res_out1 dac_3v_column_odd_0[4].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X573 dac_3v_column_0[4].dum1_in dac_3v_column_0[4].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X574 a_29905_n14015# a_31412_n14015# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X575 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X576 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X577 a_29905_n12950# dac_3v_8bit_0/b0a dac_3v_column_odd_0[4].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X578 dac_3v_8bit_0/b6a dac_3v_8bit_0/b6b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=8.4e+11p pd=8.24e+06u as=0p ps=0u w=750000u l=500000u
X579 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X580 dac_3v_8bit_0/out_unbuf dac_3v_8bit_0/b7b dac_3v_column_odd_0[6].in_5 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X581 dac_3v_column_0[4].res1_in a_22563_n12556# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X582 a_29905_n10818# dac_3v_8bit_0/b0b dac_3v_column_odd_0[3].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X583 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X584 dvdd a_n54713_n20729# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._07_.X dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X585 a_27636_2837# a_27058_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=1e+06u
X586 bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X587 a_31605_n14688# dac_3v_column_odd_0[5].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X588 dac_3v_column_odd_0[1].out1_0_3 dac_3v_8bit_0/b0a a_31605_n7227# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X589 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=8.12e+12p pd=6.412e+07u as=0p ps=0u w=2e+06u l=4e+06u
X590 dvdd in[0] a_n55547_n16609# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X591 dvss a_27998_3404# a_27636_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X592 vss follower_amp_0.nbias follower_amp_0.nbias vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X593 dvss bias_0.bi__amplifier_0.bias a_n47950_6120# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X594 testbuffer_0.tb__mux_0.tbm__passgate_1.en a_n54221_n17179# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X595 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X596 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X597 vdd level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b0b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X598 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 dvdd sky130_fd_pr__pfet_01v8_lvt ad=6.96e+12p pd=5.496e+07u as=0p ps=0u w=2e+06u l=4e+06u
X599 a_32520_2837# a_32882_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X600 a_29905_n5487# dac_3v_8bit_0/b0b dac_3v_column_0[1].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X601 a_20156_n3631# vss dac_3v_column_0[0].dum1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
D3 vss ena sky130_fd_pr__diode_pw2nd_05v5
X602 a_23802_2371# a_23802_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X603 a_33719_n16423# vdd dac_3v_column_odd_0[6].res_in0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X604 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X605 level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=4.2e+11p pd=4.12e+06u as=0p ps=0u w=750000u l=500000u
X606 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X607 dac_3v_column_odd_0[1].out1_0_0 dac_3v_8bit_0/b0a a_22563_n7227# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X608 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X609 vdd level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b0b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X610 dac_3v_column_odd_0[4].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_odd_0[4].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X611 a_20156_n13226# vdd dac_3v_column_odd_0[4].dum_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X612 testbuffer_0.tb__mux_0.tbm__passgate_4.en a_n55233_n20443# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X613 dac_3v_8bit_0/b3b dac_3v_8bit_0/b3a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X614 a_34426_n15516# vss a_34426_n15516# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X615 a_25384_n14015# dac_3v_8bit_0/b0a dac_3v_column_0[5].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X616 dac_3v_column_odd_0[4].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[4].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X617 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X618 dac_3v_column_0[5].res1_in vss a_20863_n14449# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X619 a_31942_3107# b1 dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X620 a_31412_n16147# dac_3v_8bit_0/b0b dac_3v_column_0[6].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X621 dvss dvss bandgap_0.bg__pnp_group_0.eg sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=1
X622 a_n54328_n21689# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n54400_n21689# dvss sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X623 a_33719_n2566# vss a_33719_n2566# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X624 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X625 testbuffer_0.tb__mux_0.tbm__passgate_3.en a_n54301_n18241# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X626 dvdd a_n53523_n22049# testbuffer_0.tb__mux_0.tbm__passgate_5.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X627 vdd level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=7.12e+06u w=1.5e+06u l=500000u
X628 a_25384_n7619# a_26891_n7619# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X629 dac_3v_column_0[7].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_0[7].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X630 dac_3v_column_0[5].out1_0_0 dac_3v_8bit_0/b0a a_22563_n14688# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X631 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X632 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X633 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X634 dac_3v_column_0[5].out_3 dac_3v_8bit_0/b3a dac_3v_column_0[5].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X635 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X636 dac_3v_column_odd_0[0].dum_out1 vdd a_34426_n5921# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X637 dac_3v_column_odd_0[4].out_5 dac_3v_8bit_0/b5b dac_3v_column_odd_0[4].out4 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X638 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X639 dac_3v_8bit_0/b0a dac_3v_8bit_0/b0b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=8.4e+11p pd=8.24e+06u as=0p ps=0u w=750000u l=500000u
X640 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X641 dac_3v_column_odd_0[0].res_in0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[0].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X642 dac_3v_column_0[6].out0_2 dac_3v_8bit_0/b3b dac_3v_column_0[6].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X643 dac_3v_column_0[4].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_0[4].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X644 dvss dac_3v_8bit_0/b3a dac_3v_8bit_0/b3b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X645 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.885e+13p ps=1.4334e+08u w=1e+06u l=1e+06u
X646 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X647 a_31412_n20410# vdd a_31412_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X648 dac_3v_column_0[6].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[6].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X649 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output6.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X650 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n55353_n19355# dvss dvss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X651 a_33719_n4698# vdd a_33719_n4698# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X652 dac_3v_column_odd_0[0].dum_in1 dac_3v_column_odd_0[0].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X653 a_25384_n5487# dac_3v_8bit_0/b0a dac_3v_column_0[1].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X654 a_28398_n18279# dac_3v_8bit_0/b0b dac_3v_column_0[7].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X655 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X656 a_31942_2206# a_31942_2371# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X657 vdd a_17355_n7576# vss sky130_fd_pr__res_xhigh_po w=350000u l=2.5e+07u
X658 a_33719_n11094# vss a_33719_n11094# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X659 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X660 sbamuxm4_0/ibn[0] bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[0] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X661 a_23877_n4422# dac_3v_8bit_0/b0b dac_3v_column_odd_0[0].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X662 a_25577_n17887# a_27084_n17887# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X663 a_26891_n8686# dac_3v_8bit_0/b0b dac_3v_column_odd_0[2].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X664 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X665 dac_3v_column_odd_0[4].res_out1 dac_3v_8bit_0/b0a dac_3v_column_0[5].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X666 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X667 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X668 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X669 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X670 dac_3v_column_0[0].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[0].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X671 a_23170_n4422# dac_3v_8bit_0/b2b dac_3v_column_odd_0[0].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X672 dac_3v_column_0[3].out1_0_3 dac_3v_8bit_0/b0b a_31605_n10424# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X673 dac_3v_column_odd_0[2].out0_2 dac_3v_8bit_0/b3a dac_3v_column_odd_0[2].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X674 a_32212_n2566# vss a_31605_n2963# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X675 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X676 a_29198_n2566# vss a_29198_n2566# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X677 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X678 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X679 a_n54945_n21255# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n54691_n21255# dvdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=0p ps=0u w=1e+06u l=150000u
X680 dvss level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.1e+11p ps=2.06e+06u w=750000u l=500000u
X681 dac_3v_8bit_0/b2b dac_3v_8bit_0/b2a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X682 bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inn a_n27789_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X683 dvdd a_n54301_n18241# testbuffer_0.tb__mux_0.tbm__passgate_3.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X684 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X685 dac_3v_column_odd_0[3].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_odd_0[3].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X686 a_25577_n5095# a_27084_n5095# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X687 dac_3v_column_0[5].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[5].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X688 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X689 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X690 dac_3v_column_odd_0[4].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[4].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X691 dvss a_n32029_6716# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X692 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X693 a_n54221_n16635# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output4.A dvss dvss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X694 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X695 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X696 dac_3v_8bit_0/b4a level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X697 a_25384_n19346# dac_3v_8bit_0/b0b dac_3v_column_odd_0[7].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X698 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X699 dac_3v_8bit_0/b5b dac_3v_8bit_0/b5a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X700 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X701 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X702 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X703 dvss dac_3v_8bit_0/b4a dac_3v_8bit_0/b4b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X704 a_28398_n9751# dac_3v_8bit_0/b0b dac_3v_column_0[3].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X705 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X706 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X707 dvss dac_3v_8bit_0/b5a dac_3v_8bit_0/b5b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X708 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X709 dac_3v_column_odd_0[3].out1_0_2 dac_3v_8bit_0/b0b a_27084_n11491# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X710 dvss a_33570_3107# a_34510_3404# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X711 dac_3v_column_0[0].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[0].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X712 dac_3v_column_odd_0[0].out0_2 dac_3v_8bit_0/b3b dac_3v_column_odd_0[0].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X713 dac_3v_column_odd_0[5].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[5].res_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X714 bias_0.bi__pmirr_0.gate bias_0.bi__amplifier_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=6.32e+06u as=0p ps=0u w=500000u l=1e+07u
X715 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X716 dvdd bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X717 a_34426_n9120# vss a_34426_n9120# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X718 dvss bias_0.bi__pmirr_0.gate_cas dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X719 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X720 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X721 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X722 dac_3v_column_0[0].out_3 dac_3v_8bit_0/b3b dac_3v_column_0[0].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X723 dac_3v_column_odd_0[7].out0_2 dac_3v_8bit_0/b3a dac_3v_column_odd_0[7].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X724 testbuffer_0.tb__mux_0.tbm__passgate_2.en a_n53197_n19329# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X725 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X726 a_33719_n16423# vss dac_3v_column_odd_0[6].res_in0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X727 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X728 a_23877_n18279# dac_3v_8bit_0/b0b dac_3v_column_0[7].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X729 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X730 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X731 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X732 dac_3v_8bit_0/b1a level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=8.4e+11p pd=8.24e+06u as=0p ps=0u w=750000u l=500000u
X733 dac_3v_column_0[0].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[0].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X734 dac_3v_column_0[0].out1_0_2 dac_3v_8bit_0/b0b a_27084_n4028# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X735 a_28591_n9359# a_30098_n9359# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X736 sbamuxm4_0/vb[6] a_n32029_7560# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X737 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X738 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._19_.X a_n53197_n22593# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X739 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X740 a_26891_n7619# dac_3v_8bit_0/b0a dac_3v_column_0[2].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X741 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X742 a_29905_n10818# a_31412_n10818# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X743 dac_3v_column_odd_0[2].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_odd_0[2].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X744 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X745 dac_3v_column_odd_0[7].res_in1 a_22563_n20019# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X746 a_31412_n9751# dac_3v_8bit_0/b0b dac_3v_column_0[3].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X747 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.X a_n54945_n17689# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X748 testbuffer_0.tb__mux_0.tbm__passgate_4.en a_n55233_n20443# dvss dvss sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X749 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n54945_n21255# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X750 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X751 testbuffer_0.tb__mux_0.tbm__passgate_1.en a_n54221_n17179# dvss dvss sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X752 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X753 a_20863_n2290# a_22563_n2963# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X754 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X755 a_31605_n11491# dac_3v_column_odd_0[3].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X756 sbamuxm4_0/ibn[1] bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[1] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X757 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X758 dac_3v_column_odd_0[6].out1_0_1 dac_3v_8bit_0/b0b a_24070_n17887# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X759 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X760 a_24380_2837# a_23802_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=1e+06u
X761 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n55547_n19873# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X762 dac_3v_column_odd_0[6].out_5 dac_3v_8bit_0/b5b dac_3v_column_odd_0[7].out4 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X763 a_34426_n14449# vdd a_34426_n14449# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X764 a_n40589_11895# bias_0.bi__pmirr_0.gate sbamuxm4_0/ibp[0] dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=2e+06u
X765 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X766 dac_3v_column_odd_0[6].res_in1 a_22370_n17214# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X767 a_20863_n11252# vdd a_20863_n11252# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X768 dac_3v_column_odd_0[4].out1_0_0 dac_3v_8bit_0/b0b a_22563_n13623# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X769 a_22370_n9751# dac_3v_8bit_0/b0b dac_3v_column_0[3].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X770 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X771 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X772 a_20156_n14291# vss a_20156_n14291# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X773 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X774 vdd level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=7.12e+06u w=1.5e+06u l=500000u
X775 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X776 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X777 a_n54035_n19757# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X778 dac_3v_column_odd_0[0].res_in0 dac_3v_column_odd_0[0].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X779 a_34426_n5921# vss a_34426_n5921# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X780 dac_3v_column_odd_0[7].res_in1 vdd a_20863_n19780# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X781 a_31412_n12950# dac_3v_8bit_0/b0a dac_3v_column_odd_0[4].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X782 a_31605_n9359# dac_3v_column_odd_0[2].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X783 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X784 a_30892_2837# a_31254_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X785 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X786 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X787 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X788 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X789 dac_3v_column_odd_0[2].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[2].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X790 dac_3v_column_0[2].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[2].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X791 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X792 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X793 a_n55353_n19355# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X794 level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=2.1e+11p pd=2.06e+06u as=0p ps=0u w=750000u l=500000u
X795 dac_3v_column_0[5].out1_0_1 dac_3v_8bit_0/b0b a_25577_n14688# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X796 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X797 dac_3v_column_0[1].res1_in a_22563_n6160# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X798 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbn dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X799 dac_3v_8bit_0/b7b level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X800 dvss a_31254_3404# a_30892_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X801 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X802 dac_3v_column_0[1].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_0[1].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X803 dac_3v_column_0[3].out1_0_2 dac_3v_8bit_0/b0a a_28591_n10424# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X804 a_22563_n9359# a_24070_n9359# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X805 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n48623_n18263# inp[2] dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X806 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X807 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X808 a_20156_n5763# vss a_20156_n5763# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X809 dac_3v_8bit_0/b2b dac_3v_8bit_0/b2a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X810 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X811 a_33719_n18555# vdd a_33719_n18555# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X812 follower_amp_0.vcomp dac_3v_8bit_0/out_unbuf follower_amp_0.ndrv vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X813 dac_3v_column_odd_0[2].out_5 dac_3v_8bit_0/b6b dac_3v_column_odd_0[2].in_5 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X814 dac_3v_column_0[2].out1_0_3 dac_3v_8bit_0/b0b a_30098_n8292# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X815 follower_amp_0.vcomp follower_amp_0.pbias vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X816 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X817 dac_3v_column_odd_0[3].out4 dac_3v_8bit_0/b4b dac_3v_column_odd_0[3].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X818 a_27084_n10424# a_28591_n10424# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X819 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X820 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X821 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X822 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X823 a_20863_n8053# vdd a_20863_n8053# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X824 a_22370_n17214# dac_3v_8bit_0/b0a dac_3v_column_odd_0[6].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X825 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X826 dac_3v_column_odd_0[7].res_in0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[7].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X827 dac_3v_column_0[4].out_3 dac_3v_8bit_0/b3b dac_3v_column_0[4].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X828 a_27058_3107# b4 dvss dvss sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X829 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X830 a_28398_n15082# dac_3v_8bit_0/b0b dac_3v_column_odd_0[5].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X831 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X832 dac_3v_column_0[4].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_0[4].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X833 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X834 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X835 vdd level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b7b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X836 dac_3v_column_0[2].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_0[2].res1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X837 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+12p ps=2.406e+07u w=1e+06u l=1e+06u
X838 dac_3v_column_0[1].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[1].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X839 a_33570_2371# a_34148_2837# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.142e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=1e+06u
X840 dac_3v_column_odd_0[3].res_in0 dac_3v_column_odd_0[3].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X841 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X842 dac_3v_column_odd_0[3].out1_0_3 dac_3v_8bit_0/b0b a_30098_n11491# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X843 dac_3v_column_odd_0[3].out1_0_1 dac_3v_8bit_0/b0a a_24070_n11491# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X844 dac_3v_column_odd_0[0].out1_0_1 dac_3v_8bit_0/b0a a_24070_n5095# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X845 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X846 dac_3v_8bit_0/b6b level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X847 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X848 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X849 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X850 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X851 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X852 a_23170_n19346# dac_3v_8bit_0/b2a dac_3v_column_odd_0[7].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X853 dac_3v_column_odd_0[7].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_odd_0[7].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X854 dvss a_27058_3107# a_27058_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X855 vdd level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b7b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X856 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X857 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X858 a_29905_n18279# dac_3v_8bit_0/b0b dac_3v_column_0[7].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X859 a_24070_n16820# a_25577_n16820# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X860 bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X861 dvss a_23802_3107# a_23802_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X862 level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.4e+11p pd=7.12e+06u as=0p ps=0u w=1.5e+06u l=500000u
X863 a_n42353_12343# bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=2e+06u
X864 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X865 dac_3v_8bit_0/b0b level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X866 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X867 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X868 dac_3v_8bit_0/b1b dac_3v_8bit_0/b1a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X869 dac_3v_column_0[0].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_0[0].res1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X870 a_28398_n6554# dac_3v_8bit_0/b0a dac_3v_column_odd_0[1].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X871 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X872 a_26891_n6554# a_28398_n6554# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X873 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X874 a_28591_n21083# a_30098_n21083# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X875 dac_3v_column_0[3].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_0[3].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X876 a_20156_n10027# vdd dac_3v_column_0[3].dum1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X877 a_34426_n12317# vss a_34426_n12317# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X878 dac_3v_column_0[3].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[3].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X879 testbuffer_0.tb__mux_0.tbm__passgate_3.en a_n54301_n18241# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X880 dvss level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b3a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X881 dac_3v_8bit_0/b1b dac_3v_8bit_0/b1a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X882 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X883 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X884 a_28398_n11883# dac_3v_8bit_0/b0b dac_3v_column_0[4].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X885 vdd level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b4a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X886 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X887 bias_0.bi__amplifier_0.diff bias_0.bi__amplifier_0.bias a_n47950_6120# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X888 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.32e+12p ps=1.832e+07u w=2e+06u l=1e+06u
X889 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X890 dac_3v_8bit_0/b4b dac_3v_8bit_0/b4a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X891 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X892 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X893 dvss a_28686_2206# level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X894 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X895 a_29905_n2724# vdd a_29905_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X896 a_23877_n15082# dac_3v_8bit_0/b0b dac_3v_column_odd_0[5].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X897 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X898 dac_3v_column_0[7].out1_0_1 dac_3v_8bit_0/b0a a_25577_n18952# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X899 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X900 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X901 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X902 a_29905_n4422# a_31412_n4422# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X903 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X904 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n55547_n19873# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u
X905 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n54345_n20265# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X906 a_26891_n4422# dac_3v_8bit_0/b0a dac_3v_column_odd_0[0].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X907 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X908 dac_3v_column_0[5].out1_0_3 dac_3v_8bit_0/b0b a_31605_n14688# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X909 a_31412_n6554# dac_3v_8bit_0/b0a dac_3v_column_odd_0[1].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X910 dvss a_n54443_n22593# testbuffer_0.tb__mux_0.tbm__passgate_6.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X911 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=1.032e+07u as=0p ps=0u w=1e+06u l=1e+06u
X912 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X913 a_30314_2206# a_30314_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X914 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X915 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X916 a_26184_n20686# vdd a_26184_n20686# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X917 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X918 dac_3v_column_odd_0[4].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_odd_0[4].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X919 a_n54587_n22049# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvss dvss sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X920 a_33719_n10027# vss a_33719_n10027# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X921 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X922 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X923 dvss testbuffer_0.tb__mux_0.tbm__passgate_4.en a_n47185_n21248# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X924 dvss dac_3v_8bit_0/b7b dac_3v_8bit_0/b7a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8.4e+11p ps=8.24e+06u w=750000u l=500000u
X925 dac_3v_8bit_0/out_unbuf dac_3v_8bit_0/b7a dac_3v_column_odd_0[6].in_5 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X926 a_26891_n5487# dac_3v_8bit_0/b0b dac_3v_column_0[1].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X927 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X928 a_25577_n14688# a_27084_n14688# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X929 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X930 a_33719_n18555# vss a_33719_n18555# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X931 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X932 a_23877_n9751# a_25384_n9751# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X933 a_n32750_455# dvss bandgap_0.bg__pnp_group_0.eg dvss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=9.28e+12p ps=7.328e+07u w=2e+06u l=500000u
X934 a_34426_n2724# vdd a_34426_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X935 vdd a_14987_n11444# a_14987_n11444# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X936 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X937 dac_3v_column_odd_0[6].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[6].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X938 dvss testbuffer_0.tb__mux_0.tbm__passgate_3.en a_n48623_n18263# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X939 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X940 dac_3v_column_0[1].out0_2 dac_3v_8bit_0/b3a dac_3v_column_0[1].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X941 a_30098_n18952# a_31605_n18952# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X942 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X943 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inp bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.64e+12p ps=3.432e+07u w=4e+06u l=1e+06u
X944 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X945 vdd dac_3v_8bit_0/b7b dac_3v_8bit_0/b7a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X946 dac_3v_column_odd_0[7].out1_0_0 dac_3v_8bit_0/b0a a_22563_n20019# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X947 dac_3v_column_odd_0[4].out1_0_2 dac_3v_8bit_0/b0a a_27084_n13623# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X948 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X949 dvss a_n55547_n19873# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X950 a_23170_n4422# dac_3v_8bit_0/b1a dac_3v_column_odd_0[0].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X951 dac_3v_column_odd_0[7].out_3 dac_3v_8bit_0/b3a dac_3v_column_odd_0[7].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X952 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output5.A a_n54035_n19757# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X953 a_30705_n2566# vdd a_30705_n2566# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X954 a_20024_n21083# a_20863_n20410# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X955 dac_3v_column_odd_0[2].res_in0 dac_3v_column_odd_0[2].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X956 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbn dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X957 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X958 a_23877_n11883# dac_3v_8bit_0/b0b dac_3v_column_0[4].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X959 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X960 dac_3v_column_odd_0[2].out1_0_3 dac_3v_8bit_0/b0a a_30098_n9359# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X961 dac_3v_column_0[2].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[2].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X962 dvss bias_0.bi__nmirr_0.gate_n a_n42000_7938# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X963 a_20863_n2290# vdd a_20863_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X964 a_25384_n2724# vdd a_25384_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X965 a_28591_n2963# a_30098_n2963# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X966 dac_3v_column_odd_0[5].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_odd_0[5].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X967 a_n46909_n21248# a_n47185_n21248# dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X968 dvss testbuffer_0.tb__mux_0.tbm__passgate_6.en a_n47185_n24233# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X969 dac_3v_column_odd_0[3].out1_0_3 dac_3v_8bit_0/b0a a_30098_n11491# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X970 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X971 dvdd a_n54443_n22593# testbuffer_0.tb__mux_0.tbm__passgate_6.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X972 a_25384_n16147# dac_3v_8bit_0/b0b dac_3v_column_0[6].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X973 a_n32750_n2725# dvss bandgap_0.bg__pnp_group_0.eg dvss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X974 dvdd in[1] a_n55547_n19873# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X975 a_23877_n20410# a_25384_n20410# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X976 a_n21613_n925# a_n21227_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X977 dvss a_n55547_n16609# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X978 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output6.A a_n55047_n18669# a_n54937_n18785# dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X979 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C a_n54328_n21689# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X980 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X981 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output4.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X982 dac_3v_column_odd_0[2].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[2].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X983 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X984 a_21663_n2566# vdd a_21663_n2566# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X985 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X986 a_22563_n15755# a_24070_n15755# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X987 dac_3v_column_odd_0[7].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_odd_0[7].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X988 a_33719_n15358# vdd a_33719_n15358# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X989 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X990 level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=4.2e+11p pd=4.12e+06u as=0p ps=0u w=750000u l=500000u
X991 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X992 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X993 dac_3v_column_0[7].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_0[7].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X994 dac_3v_column_0[4].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_0[4].res1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X995 dvdd a_n53983_n17697# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X996 a_20863_n18713# vss a_20863_n18713# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X997 dac_3v_column_odd_0[4].out_5 dac_3v_8bit_0/b5a dac_3v_column_odd_0[4].out4 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X998 dac_3v_8bit_0/b5a level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X999 dac_3v_column_0[3].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[3].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1000 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1001 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out a_n23132_n3629# dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X1002 dac_3v_column_0[6].out0_2 dac_3v_8bit_0/b3a dac_3v_column_0[6].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1003 a_26891_n15082# a_28398_n15082# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1004 dvdd bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=1.264e+07u w=500000u l=2e+06u
X1005 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1006 a_n54713_n20729# a_n54440_n20729# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.5725e+11p pd=2.99e+06u as=0p ps=0u w=420000u l=150000u
X1007 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1008 a_n32750_n4845# dvss bandgap_0.bg__pnp_group_0.eg dvss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1009 a_25384_n20410# vdd a_25384_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1010 dvdd bias_0.bi__amplifier_0.mirr bias_0.bi__pmirr_0.gate dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X1011 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1012 a_n48347_n18263# a_n48623_n18263# dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1013 a_31605_n2963# vhigh vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1014 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1015 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1016 a_20863_n20410# vss a_20863_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1017 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.A a_n54945_n17689# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1018 vdd follower_amp_0.pbias follower_amp_0.pbias vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1019 a_28591_n6160# a_30098_n6160# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1020 dac_3v_column_odd_0[2].res_in1 vss a_20863_n9120# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1021 a_24070_n7227# a_25577_n7227# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1022 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1023 dac_3v_8bit_0/b3a level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1024 a_26891_n17214# dac_3v_8bit_0/b0b dac_3v_column_odd_0[6].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1025 dac_3v_column_odd_0[2].res_in0 dac_3v_column_odd_0[2].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1026 dac_3v_column_odd_0[1].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_odd_0[1].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1027 dvss a_22174_3107# a_23114_3404# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X1028 dac_3v_8bit_0/b0a dac_3v_8bit_0/b0b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1029 a_22370_n17214# dac_3v_8bit_0/b0b dac_3v_column_odd_0[6].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1030 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n54072_n20437# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.087e+11p ps=1.36e+06u w=420000u l=150000u
X1031 dac_3v_column_odd_0[0].out4 dac_3v_8bit_0/b4a dac_3v_column_odd_0[0].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1032 a_23170_n20686# vdd a_22563_n21083# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1033 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1034 dvss level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1035 dac_3v_column_0[1].out1_0_3 dac_3v_8bit_0/b0a a_30098_n6160# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1036 a_26891_n20844# vss a_26891_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1037 dac_3v_column_odd_0[5].res_in0 dac_3v_column_odd_0[5].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1038 dvss bias_0.bi__nmirr_0.gate_n dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1039 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1040 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._19_.X a_n53289_n21505# dvss dvss sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1041 a_23170_n6554# dac_3v_8bit_0/b1a dac_3v_column_odd_0[1].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1042 dac_3v_8bit_0/b7b level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1043 a_22563_n2963# a_24070_n2963# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1044 dac_3v_column_odd_0[2].out1_0_1 dac_3v_8bit_0/b0b a_25577_n9359# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1045 a_n53615_n20961# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1046 a_29905_n15082# dac_3v_8bit_0/b0b dac_3v_column_odd_0[5].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1047 a_24070_n13623# a_25577_n13623# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1048 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1049 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1050 dac_3v_column_0[5].res1_in a_22370_n14015# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1051 dac_3v_column_0[1].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_0[1].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1052 a_n55547_n16609# in[0] dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1053 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1054 dac_3v_column_0[5].out1_0_2 dac_3v_8bit_0/b0a a_28591_n14688# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1055 dac_3v_column_0[3].out1_0_0 dac_3v_8bit_0/b0b a_22563_n10424# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1056 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1057 a_27058_2206# a_27058_2371# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X1058 dvss a_31254_3404# a_30892_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1059 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output4.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1060 dac_3v_column_odd_0[7].out4 dac_3v_8bit_0/b4b dac_3v_column_0[7].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1061 dac_3v_column_odd_0[5].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[5].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1062 a_33719_n12159# vdd a_33719_n12159# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1063 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1064 dac_3v_column_odd_0[0].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[0].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1065 dvss level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4.2e+11p ps=4.12e+06u w=750000u l=500000u
X1066 a_31605_n6160# dac_3v_column_odd_0[1].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1067 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1068 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1069 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1070 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1071 dac_3v_column_0[6].res1_in vdd a_20863_n16581# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1072 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1073 a_n54221_n16635# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output4.A dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1074 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1075 dac_3v_column_odd_0[1].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_odd_0[1].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1076 a_23170_n12950# dac_3v_8bit_0/b1a dac_3v_column_odd_0[4].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1077 a_20156_n8962# vdd a_20156_n8962# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1078 dac_3v_column_0[2].out1_0_2 dac_3v_8bit_0/b0a a_28591_n8292# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1079 dvss bias_0.bi__nmirr_0.gate_n a_n42000_7586# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1080 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1081 vlow vss a_32919_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1082 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1083 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1084 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1085 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1086 vdd dac_3v_8bit_0/b3a dac_3v_8bit_0/b3b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1087 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1088 level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.4e+11p pd=7.12e+06u as=0p ps=0u w=1.5e+06u l=500000u
X1089 dac_3v_column_0[7].out1_0_2 dac_3v_8bit_0/b0b a_28591_n18952# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1090 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n55353_n19355# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1091 dac_3v_column_odd_0[6].dum_in0 vss a_34426_n17648# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1092 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1093 a_22563_n6160# a_24070_n6160# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1094 dac_3v_column_odd_0[6].out1_0_3 dac_3v_8bit_0/b0a a_31605_n17887# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1095 dac_3v_column_odd_0[5].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[5].res_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X1096 a_20863_n3789# vss a_20863_n3789# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1097 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1098 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C a_n54440_n20729# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.087e+11p ps=1.36e+06u w=420000u l=150000u
X1099 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1100 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1101 a_34426_n19780# vdd a_34426_n19780# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1102 a_29198_n20686# vss a_29198_n20686# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1103 a_n54195_n20411# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C dvss dvss sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=0p ps=0u w=420000u l=150000u
X1104 dac_3v_8bit_0/b1a level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1105 dac_3v_column_odd_0[0].out_5 dac_3v_8bit_0/b5a dac_3v_column_odd_0[1].out4 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1106 dac_3v_column_0[1].out1_0_1 dac_3v_8bit_0/b0b a_25577_n6160# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1107 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1108 dac_3v_8bit_0/b7b level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1109 a_29905_n11883# dac_3v_8bit_0/b0b dac_3v_column_0[4].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1110 dac_3v_column_0[2].out1_0_3 dac_3v_8bit_0/b0a a_31605_n8292# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1111 vdd level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1112 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1113 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1114 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1115 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1116 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1117 dac_3v_column_odd_0[5].res_out1 dac_3v_8bit_0/b0b dac_3v_column_0[6].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1118 a_22370_n14015# dac_3v_8bit_0/b0a dac_3v_column_0[5].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1119 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.64e+12p ps=3.432e+07u w=4e+06u l=1e+06u
X1120 testbuffer_0.tb__mux_0.tbm__passgate_6.en a_n54443_n22593# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1121 a_22174_2371# a_22752_2837# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.142e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=1e+06u
X1122 a_29905_n19346# a_31412_n19346# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1123 dac_3v_8bit_0/b1a level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1124 dac_3v_column_odd_0[7].out1_0_1 dac_3v_8bit_0/b0b a_25577_n20019# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1125 a_33719_n15358# vss a_33719_n15358# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1126 a_25577_n11491# a_27084_n11491# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1127 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1128 dac_3v_column_0[2].out1_0_0 dac_3v_8bit_0/b0a a_22563_n8292# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1129 a_20156_n3631# vdd dac_3v_column_0[0].dum1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1130 dac_3v_column_0[5].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_0[5].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1131 a_20156_n14291# vdd dac_3v_column_0[5].dum1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1132 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1133 a_20156_n2566# vss a_20024_n2963# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1134 dac_3v_column_0[5].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[5].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1135 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1136 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1137 a_28686_2206# a_28686_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X1138 a_33719_n15358# vdd dac_3v_column_odd_0[5].res_out1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1139 bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1140 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1141 dac_3v_column_0[6].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_0[6].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1142 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1143 dac_3v_column_0[6].out0_1_1 dac_3v_8bit_0/b2a dac_3v_column_0[6].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1144 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inn bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1145 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n48623_n21248# inp[5] dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1146 a_33570_2371# a_33570_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X1147 dac_3v_8bit_0/b4b dac_3v_8bit_0/b4a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1148 a_22370_n18279# a_23877_n18279# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1149 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1150 a_25384_n12950# dac_3v_8bit_0/b0a dac_3v_column_odd_0[4].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1151 a_n53553_n18785# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n53825_n18785# dvdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=0p ps=0u w=1e+06u l=150000u
X1152 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1153 dac_3v_column_odd_0[0].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[0].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1154 dac_3v_column_odd_0[4].res_in1 vss a_20863_n13384# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1155 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1156 a_13761_n11418# dac_out follower_amp_0.vcomp vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X1157 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1158 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n55547_n19873# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1159 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1160 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1161 a_20156_n18555# vss dac_3v_column_0[7].dum1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1162 vdd level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b2a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1163 a_28398_n3355# dac_3v_8bit_0/b0a dac_3v_column_0[0].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1164 a_34426_n20844# vdd a_34426_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1165 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1166 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1167 a_26891_n3355# a_28398_n3355# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1168 dac_3v_column_odd_0[6].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_odd_0[6].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1169 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1170 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1171 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n53983_n17697# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1172 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1173 a_23170_n10818# dac_3v_8bit_0/b1b dac_3v_column_odd_0[3].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1174 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1175 testbuffer_0.tb__mux_0.tbm__passgate_6.en a_n54443_n22593# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1176 dvss a_28686_3107# a_28686_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1177 a_26891_n10818# dac_3v_8bit_0/b0a dac_3v_column_odd_0[3].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1178 vdd a_27058_2206# level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X1179 a_20156_n20686# vss a_20156_n20686# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1180 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1181 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1182 dac_3v_column_odd_0[1].out1_0_0 dac_3v_8bit_0/b0b a_22563_n7227# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1183 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1184 a_29905_n16147# a_31412_n16147# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1185 level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1186 vdd follower_amp_0.pbias follower_amp_0.vcomp vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1187 dvss bias_0.bi__amplifier_0.bias bias_0.bi__amplifier_0.bias dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=1.264e+07u w=500000u l=4e+06u
X1188 dac_3v_column_odd_0[5].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[5].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1189 a_33719_n12159# vss a_33719_n12159# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1190 dac_3v_column_odd_0[6].out_5 dac_3v_8bit_0/b6b dac_3v_column_odd_0[6].in_5 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1191 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1192 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inn bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1193 a_n53983_n17697# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1194 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1195 a_31605_n16820# dac_3v_column_odd_0[6].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1196 a_26184_n20686# vss a_25577_n21083# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1197 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1198 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1199 a_31412_n3355# dac_3v_8bit_0/b0a dac_3v_column_0[0].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1200 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1201 dac_3v_column_odd_0[4].res_in0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[4].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1202 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1203 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1204 a_29905_n7619# dac_3v_8bit_0/b0b dac_3v_column_0[2].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1205 bias_0.bi__nmirr_0.gate_n bias_0.bi__nmirr_0.gate_n dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=1.032e+07u as=0p ps=0u w=1e+06u l=2e+06u
X1206 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1207 dac_3v_8bit_0/b1a level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1208 a_29198_n2566# vdd a_29198_n2566# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1209 dac_3v_column_odd_0[3].out1_0_1 dac_3v_8bit_0/b0b a_24070_n11491# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1210 dac_3v_column_0[3].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_0[3].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1211 a_n32750_n605# dvdd bandgap_0.bg__pnp_group_0.eg dvss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1212 dac_3v_column_odd_0[3].res_in1 a_22370_n10818# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1213 a_n54221_n17179# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output5.A dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1214 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1215 vdd level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b3a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1216 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1217 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1218 a_27058_2371# a_27636_2837# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.142e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=1e+06u
X1219 a_23170_n19346# dac_3v_8bit_0/b2b dac_3v_column_odd_0[7].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1220 dac_3v_column_odd_0[4].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[4].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1221 a_n32750_n605# a_n31275_n1537# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1222 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1223 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1224 a_25384_n9751# a_26891_n9751# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1225 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1226 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1227 dac_3v_column_0[6].out1_0_0 dac_3v_8bit_0/b0a a_22563_n16820# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1228 dac_3v_column_0[3].out1_0_2 dac_3v_8bit_0/b0a a_27084_n10424# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1229 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1230 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n54657_n18785# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1231 a_n55233_n20443# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output8.A dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1232 dac_3v_8bit_0/b7a dac_3v_8bit_0/b7b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1233 a_28398_n8686# dac_3v_8bit_0/b0b dac_3v_column_odd_0[2].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1234 a_n42353_11447# bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=2e+06u
X1235 dac_3v_column_0[6].out_3 dac_3v_8bit_0/b3a dac_3v_column_0[6].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1236 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1237 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1238 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1239 dac_3v_8bit_0/b5b dac_3v_8bit_0/b5a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1240 dac_3v_column_odd_0[0].res_out1 dac_3v_column_odd_0[0].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1241 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1242 dac_3v_column_odd_0[1].dum_out1 vdd a_34426_n8053# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1243 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1244 dvdd a_n53523_n22049# testbuffer_0.tb__mux_0.tbm__passgate_5.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1245 dac_3v_column_odd_0[2].out4 dac_3v_8bit_0/b4b dac_3v_column_odd_0[2].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1246 a_32212_n2566# vdd a_32212_n2566# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1247 dac_3v_column_odd_0[7].out1_0_3 dac_3v_8bit_0/b0b a_31605_n20019# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1248 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1249 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1250 a_n32750_n2725# a_n31275_n3657# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1251 dac_3v_column_0[4].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_0[4].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1252 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1253 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1254 a_33719_n8962# vdd dac_3v_column_odd_0[2].res_out1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X1255 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1256 a_26891_n2724# vdd a_26891_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1257 a_33719_n15358# vss dac_3v_column_odd_0[5].res_out1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X1258 bias_0.bi__amplifier_0.bias bias_0.bi__amplifier_0.bias dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1259 dvdd a_27058_3107# a_27998_3404# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X1260 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1261 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1262 dac_3v_column_odd_0[1].dum_in1 dac_3v_column_odd_0[1].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1263 a_22563_n12556# a_24070_n12556# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1264 a_25384_n7619# dac_3v_8bit_0/b0a dac_3v_column_0[2].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1265 dac_3v_column_0[6].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_0[6].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1266 dac_3v_column_odd_0[2].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[2].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1267 dvss level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b2a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1268 a_23170_n2566# vdd a_23170_n2566# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1269 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1270 a_27691_n2566# vdd a_27084_n2963# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1271 dvdd bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1272 a_31412_n8686# dac_3v_8bit_0/b0b dac_3v_column_odd_0[2].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X1273 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1274 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1275 dac_3v_column_odd_0[2].out1_0_1 dac_3v_8bit_0/b0b a_24070_n9359# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1276 a_n32750_n4845# bandgap_0.bg__pnp_group_0.eg dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1277 a_26891_n11883# a_28398_n11883# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1278 dac_3v_column_0[3].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_0[3].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1279 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1280 a_33570_3107# b0 dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X1281 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1282 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1283 dac_3v_column_0[5].out1_0_0 dac_3v_8bit_0/b0b a_22563_n14688# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1284 dvdd bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1285 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inp bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1286 vdd level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1287 dac_3v_column_0[3].res1_in vdd a_20863_n10185# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1288 bias_0.bi__nmirr_0.gate_n bias_0.bi__nmirr_0.gate_n dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1289 a_30314_3107# b2 dvss dvss sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X1290 a_24070_n4028# a_25577_n4028# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1291 dac_3v_column_0[1].res1_in vss a_20863_n5921# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1292 a_26891_n14015# dac_3v_8bit_0/b0b dac_3v_column_0[5].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1293 dac_3v_column_odd_0[4].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_odd_0[4].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1294 dac_3v_column_odd_0[3].dum_in0 vdd a_34426_n11252# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1295 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1296 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1297 a_22370_n8686# dac_3v_8bit_0/b0b dac_3v_column_odd_0[2].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1298 a_25577_n7227# a_27084_n7227# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1299 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1300 dac_3v_column_0[0].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_0[0].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1301 dac_3v_column_odd_0[1].out4 dac_3v_8bit_0/b4a dac_3v_column_0[1].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1302 a_22370_n14015# dac_3v_8bit_0/b0b dac_3v_column_0[5].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1303 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1304 a_20156_n13226# vss a_20156_n13226# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1305 dvss a_n53197_n19329# testbuffer_0.tb__mux_0.tbm__passgate_2.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1306 testbuffer_0.tb__mux_0.tbm__passgate_5.en a_n53523_n22049# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1307 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1308 a_31412_n20410# vlow vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1309 dac_3v_column_odd_0[2].out_5 dac_3v_8bit_0/b5b dac_3v_column_odd_0[3].out4 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1310 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1311 dac_3v_column_odd_0[3].res_out1 dac_3v_column_odd_0[3].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1312 dac_3v_column_0[0].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[0].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1313 a_34426_n4856# vss a_34426_n4856# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1314 dac_3v_8bit_0/b0a dac_3v_8bit_0/b0b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1315 vdd dac_3v_8bit_0/b4a dac_3v_8bit_0/b4b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1316 a_33719_n5763# vdd dac_3v_column_odd_0[1].res_in0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X1317 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1318 vdd level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b1a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1319 a_24070_n10424# a_25577_n10424# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1320 a_23170_n6554# dac_3v_8bit_0/b2a dac_3v_column_odd_0[1].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1321 testbuffer_0.tb__mux_0.tbm__passgate_0.en a_n54221_n16635# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1322 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n48347_n21248# inp[5] dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1323 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1324 a_32212_n20686# vss a_31605_n21083# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1325 dac_3v_column_odd_0[2].out1_0_2 dac_3v_8bit_0/b0a a_27084_n9359# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1326 dac_3v_column_odd_0[4].out1_0_2 dac_3v_8bit_0/b0b a_27084_n13623# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1327 dvss a_30314_3107# a_30314_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1328 dac_3v_column_0[1].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[1].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1329 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1330 dac_3v_column_0[4].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[4].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1331 a_23170_n10818# dac_3v_8bit_0/b1b dac_3v_column_odd_0[3].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1332 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1333 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1334 dac_3v_8bit_0/b1a level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1335 dvss a_31942_2206# level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X1336 dac_3v_column_odd_0[0].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_odd_0[0].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1337 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1338 sbamuxm4_0/ibn[0] bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[0] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1339 a_11923_n8212# a_17355_n8212# vss sky130_fd_pr__res_xhigh_po w=350000u l=2.5e+07u
X1340 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1341 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inp bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1342 a_20156_n5763# vdd a_20156_n5763# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1343 dac_3v_column_0[0].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_0[0].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1344 dac_3v_column_0[1].out1_0_1 dac_3v_8bit_0/b0b a_24070_n6160# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1345 dvdd a_n55547_n16609# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1346 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1347 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1348 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1349 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1350 dvdd a_n54345_n20265# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.X dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1351 level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X1352 dvss level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b0b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1353 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1354 a_29905_n12950# a_31412_n12950# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1355 dac_3v_column_odd_0[4].dum_out1 vss a_34426_n14449# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1356 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1357 dac_3v_column_0[4].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_0[4].res1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X1358 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1359 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n48347_n24233# inp[6] dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1360 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1361 dvss level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1362 a_31605_n13623# dac_3v_column_odd_0[4].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1363 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1364 dac_3v_column_0[0].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_0[0].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1365 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1366 a_28686_2371# a_28686_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1367 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1368 a_34426_n16581# vdd a_34426_n16581# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1369 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1370 a_20863_n13384# vdd a_20863_n13384# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1371 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1372 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1373 dac_3v_column_odd_0[0].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[0].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1374 dac_3v_column_odd_0[7].out1_0_2 dac_3v_8bit_0/b0a a_28591_n20019# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1375 dac_3v_8bit_0/b5a level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.68e+12p pd=1.424e+07u as=0p ps=0u w=1.5e+06u l=500000u
X1376 a_29905_n4422# dac_3v_8bit_0/b0b dac_3v_column_odd_0[0].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1377 dac_3v_column_0[1].out1_0_2 dac_3v_8bit_0/b0a a_27084_n6160# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1378 dvdd bias_0.bi__amplifier_0.mirr bias_0.bi__pmirr_0.gate dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X1379 a_n54221_n17179# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output5.A dvss dvss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1380 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output8.A a_n54441_n21531# dvss dvss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X1381 dvss dac_3v_8bit_0/b5a dac_3v_8bit_0/b5b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1382 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1383 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbn dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1384 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X a_n53983_n17697# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1385 vdd level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1386 a_n46909_n15278# a_n47185_n15278# dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1387 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1388 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1389 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1390 dac_3v_column_0[6].out1_0_1 dac_3v_8bit_0/b0b a_25577_n16820# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1391 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1392 a_26891_n7619# a_28398_n7619# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1393 a_n55547_n16609# in[0] dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1394 a_28591_n15755# a_30098_n15755# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1395 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n53615_n20961# dvss dvss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X1396 dvss a_33570_3107# a_33570_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1397 a_33719_n12159# vdd dac_3v_column_odd_0[4].res_in0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1398 dac_3v_column_odd_0[3].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[3].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1399 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1400 a_21663_n2566# vss a_20863_n2290# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1401 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1402 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n55353_n19355# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1403 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1404 vdd dac_3v_8bit_0/b6b dac_3v_8bit_0/b6a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1405 dac_3v_8bit_0/b2a level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1406 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1407 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X a_n55547_n16609# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1408 a_32919_n2290# a_32919_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1409 dac_3v_column_odd_0[0].dum_in0 vdd a_34426_n4856# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1410 a_n55681_n18241# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.415e+11p pd=2.83e+06u as=0p ps=0u w=420000u l=150000u
X1411 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1412 a_20156_n7895# vss a_20156_n7895# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1413 a_29905_n19346# dac_3v_8bit_0/b0a dac_3v_column_odd_0[7].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1414 level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=2.1e+11p pd=2.06e+06u as=0p ps=0u w=750000u l=500000u
X1415 dvss dac_3v_8bit_0/b6b dac_3v_8bit_0/b6a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1416 a_n42353_12567# bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1417 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1418 dac_3v_column_odd_0[4].out4 dac_3v_8bit_0/b4b dac_3v_column_odd_0[4].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1419 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1420 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output4.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1421 a_n54487_n21933# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1422 dac_3v_column_0[7].res1_in a_22563_n18952# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1423 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output7.A a_n55313_n22049# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1424 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1425 a_22563_n20019# a_24070_n20019# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1426 dac_3v_column_odd_0[0].res_in1 a_22370_n4422# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1427 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1428 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1429 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._19_.A a_n54487_n21933# dvss dvss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1430 follower_amp_0.nbias follower_amp_0.nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1431 dvdd bias_0.bi__pmirr_0.gate a_n40589_12343# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X1432 level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1433 vdd dac_3v_8bit_0/b5a dac_3v_8bit_0/b5b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1434 a_28398_n17214# dac_3v_8bit_0/b0b dac_3v_column_odd_0[6].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X1435 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output6.A a_n54301_n18241# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1436 a_25384_n4422# dac_3v_8bit_0/b0a dac_3v_column_odd_0[0].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1437 a_29198_n20686# vdd a_28591_n21083# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1438 dac_3v_column_odd_0[6].out1_0_1 dac_3v_8bit_0/b0a a_25577_n17887# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1439 sbamuxm4_0/vb[1] a_n32029_10936# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1440 dvdd testbuffer_0.tb__mux_0.tbm__passgate_3.en a_n48623_n18263# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1441 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1442 a_22174_2371# a_22174_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X1443 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1444 dac_3v_8bit_0/b1b dac_3v_8bit_0/b1a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1445 dac_3v_column_0[7].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[7].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1446 a_22370_n17214# a_23877_n17214# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1447 dac_3v_column_0[5].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_0[5].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1448 level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1449 a_26891_n18279# dac_3v_8bit_0/b0a dac_3v_column_0[7].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1450 a_20156_n19622# vdd dac_3v_column_odd_0[7].dum_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1451 dac_3v_column_odd_0[7].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_odd_0[7].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1452 dac_3v_column_odd_0[4].out1_0_3 dac_3v_8bit_0/b0b a_30098_n13623# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1453 dac_3v_column_odd_0[4].out1_0_1 dac_3v_8bit_0/b0a a_24070_n13623# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1454 dvss level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1455 dac_3v_column_odd_0[3].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[3].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1456 dac_3v_column_odd_0[1].out1_0_1 dac_3v_8bit_0/b0a a_24070_n7227# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1457 vdd dac_3v_8bit_0/b3a dac_3v_8bit_0/b3b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1458 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1459 dac_3v_column_odd_0[7].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[7].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1460 dac_3v_column_0[4].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[4].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1461 a_n54114_n20411# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n54195_n20411# dvss sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X1462 dac_3v_column_odd_0[4].out_5 dac_3v_8bit_0/b5a dac_3v_column_odd_0[5].out4 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1463 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1464 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1465 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1466 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n54441_n21531# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1467 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1468 sbamuxm4_0/ibn[1] bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[1] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1469 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
D4 vss dac_3v_8bit_0/out_unbuf sky130_fd_pr__diode_pw2nd_05v5
X1470 a_33719_n8962# vss a_33719_n8962# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1471 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1472 dvss a_n53615_n20961# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1473 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1474 dvdd testbuffer_0.tb__mux_0.tbm__passgate_6.en a_n47185_n24233# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1475 a_27084_n5095# a_28591_n5095# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1476 dvss a_n55353_n19355# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1477 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1478 dac_3v_8bit_0/b7b level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1479 dac_3v_column_0[5].out1_0_2 dac_3v_8bit_0/b0a a_27084_n14688# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1480 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1481 a_23877_n8686# a_25384_n8686# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1482 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1483 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1484 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1485 a_30098_n17887# a_31605_n17887# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1486 dac_3v_column_odd_0[5].dum_in1 dac_3v_column_odd_0[5].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1487 dac_3v_8bit_0/b3a level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1488 dac_3v_column_0[7].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_0[7].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1489 a_n32750_n1665# dvss bandgap_0.bg__pnp_group_0.eg dvss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1490 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1491 dac_3v_column_odd_0[1].res_in0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[1].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1492 dvss bias_0.bi__pmirr_0.gate_cas dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1493 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1494 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1495 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1496 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1497 dac_3v_column_0[6].out0_1_1 dac_3v_8bit_0/b2b dac_3v_column_0[6].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1498 dvss dvss bandgap_0.bg__pnp_group_0.eg sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=1
X1499 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1500 a_23877_n15082# a_25384_n15082# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1501 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1502 a_22370_n20410# vdd a_22370_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1503 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1504 testbuffer_0.tb__mux_0.tbm__passgate_3.en a_n54301_n18241# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1505 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1506 a_30314_2206# a_30314_2371# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X1507 follower_amp_0.vcomp dac_out a_13761_n11418# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1508 dac_3v_8bit_0/b4b dac_3v_8bit_0/b4a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1509 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1510 a_28398_n5487# dac_3v_8bit_0/b0b dac_3v_column_0[1].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1511 bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1512 a_23877_n17214# dac_3v_8bit_0/b0b dac_3v_column_odd_0[6].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1513 a_23877_n6554# dac_3v_8bit_0/b0a dac_3v_column_odd_0[1].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X1514 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inp bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1515 a_n32750_n3785# dvss bandgap_0.bg__pnp_group_0.eg dvss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1516 dvss a_n54221_n16635# testbuffer_0.tb__mux_0.tbm__passgate_0.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1517 dac_3v_column_odd_0[2].out_3 dac_3v_8bit_0/b3a dac_3v_column_odd_0[2].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1518 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1519 a_29905_n6554# a_31412_n6554# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1520 dac_3v_column_odd_0[6].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_odd_0[6].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1521 a_20156_n20686# vdd a_20024_n21083# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1522 a_28398_n20844# vdd a_28398_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1523 dac_3v_8bit_0/b4b dac_3v_8bit_0/b4a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1524 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1525 dac_3v_column_0[6].out1_0_3 dac_3v_8bit_0/b0b a_31605_n16820# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1526 dac_3v_column_0[3].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[3].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1527 a_23877_n20844# vss a_23877_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1528 a_20863_n17648# vss a_20863_n17648# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1529 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.A a_n54945_n17689# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1530 a_33719_n3631# vss dac_3v_column_odd_0[0].res_in0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X1531 dac_3v_column_odd_0[2].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[2].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1532 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1533 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1534 dac_3v_column_odd_0[3].out1_0_3 dac_3v_8bit_0/b0a a_31605_n11491# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1535 a_n48347_n21248# a_n48623_n21248# dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1536 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1537 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1538 level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1539 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1540 dvss dvdd w_n19679_n3822# w_n19679_n3822# sky130_fd_pr__pfet_01v8 ad=3.44222e+14p pd=3.50579e+09u as=5.8e+11p ps=5.16e+06u w=1e+06u l=1e+06u
X1541 a_33719_n12159# vss dac_3v_column_odd_0[4].res_in0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1542 a_24070_n8292# a_25577_n8292# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1543 dac_3v_column_0[2].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_0[2].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1544 dvss a_n54443_n22593# testbuffer_0.tb__mux_0.tbm__passgate_6.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1545 dac_3v_column_0[0].dum1_in dac_3v_column_0[0].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1546 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1547 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1548 dac_3v_column_odd_0[7].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[7].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1549 dac_3v_column_odd_0[6].out_5 dac_3v_8bit_0/b6a dac_3v_column_odd_0[6].in_5 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1550 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1551 a_26891_n7619# dac_3v_8bit_0/b0b dac_3v_column_0[2].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1552 sbamuxm4_0/vb[4] a_n32029_9248# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1553 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1554 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1555 follower_amp_0.nbias ena a_11923_n8212# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1556 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1557 a_25577_n16820# a_27084_n16820# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1558 a_n53925_n19873# a_n54035_n19757# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output5.A dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1559 a_31412_n5487# dac_3v_8bit_0/b0b dac_3v_column_0[1].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X1560 a_22174_3107# b7 dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X1561 a_28398_n18279# a_29905_n18279# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1562 bias_0.bi__pmirr_0.fb bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1563 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1564 dac_3v_column_odd_0[0].out1_0_3 dac_3v_8bit_0/b0a a_30098_n5095# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1565 dac_3v_column_odd_0[2].out1_0_1 dac_3v_8bit_0/b0a a_25577_n9359# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1566 dac_3v_column_0[2].out0_2 dac_3v_8bit_0/b3a dac_3v_column_0[2].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1567 dvdd bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1568 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1569 dvss a_31942_3107# a_32882_3404# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X1570 dac_3v_8bit_0/b7b level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1571 dac_3v_column_0[3].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[3].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1572 bias_0.bi__amplifier_0.diff bias_0.bi__amplifier_0.inn bias_0.bi__pmirr_0.gate dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X1573 dvss a_n55233_n20443# testbuffer_0.tb__mux_0.tbm__passgate_4.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1574 a_n48347_n24233# a_n48623_n24233# dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1575 dvss dac_3v_8bit_0/b6b dac_3v_8bit_0/b6a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1576 dac_3v_column_0[3].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_0[3].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1577 vdd level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b5a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1578 dac_3v_column_odd_0[0].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[0].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1579 bias_0.bi__amplifier_0.bias bias_0.bi__amplifier_0.bias dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1580 a_25577_n4028# a_27084_n4028# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1581 a_22370_n5487# dac_3v_8bit_0/b0b dac_3v_column_0[1].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1582 dac_3v_column_0[1].out_3 dac_3v_8bit_0/b3a dac_3v_column_0[1].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1583 dac_3v_column_odd_0[6].out4 dac_3v_8bit_0/b4a dac_3v_column_odd_0[6].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1584 dac_3v_column_0[2].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_0[2].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1585 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1586 dvss a_n55547_n19873# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1587 dac_3v_8bit_0/b5b dac_3v_8bit_0/b5a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1588 dac_3v_column_odd_0[6].dum_out1 vdd a_34426_n18713# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1589 dac_3v_column_odd_0[3].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[3].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1590 dac_3v_8bit_0/b1a level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1591 dac_3v_column_odd_0[4].out1_0_3 dac_3v_8bit_0/b0a a_30098_n13623# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1592 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1593 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1594 dac_3v_column_0[3].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[3].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1595 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1596 dac_3v_8bit_0/b2b dac_3v_8bit_0/b2a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1597 dac_3v_column_odd_0[7].res_in1 a_22370_n19346# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1598 dvss a_31942_3107# a_31942_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1599 a_31942_2206# a_31942_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X1600 dac_3v_column_0[0].out0_1_1 dac_3v_8bit_0/b2a dac_3v_column_0[0].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1601 dac_3v_column_0[0].out1_0_2 dac_3v_8bit_0/b0b a_28591_n4028# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1602 a_20156_n4698# vss a_20156_n4698# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1603 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1604 a_33719_n17490# vdd a_33719_n17490# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1605 dvdd a_n54443_n22593# testbuffer_0.tb__mux_0.tbm__passgate_6.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1606 vdd a_30314_2206# level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X1607 dvss level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b4a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1608 dac_3v_column_0[3].out1_0_2 dac_3v_8bit_0/b0b a_27084_n10424# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1609 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1610 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1611 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1612 level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=2.1e+11p pd=2.06e+06u as=0p ps=0u w=750000u l=500000u
X1613 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1614 dac_3v_column_odd_0[6].out1_0_2 dac_3v_8bit_0/b0b a_28591_n17887# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1615 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1616 sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=3.48e+12p pd=2.574e+07u as=0p ps=0u w=4e+06u l=4e+06u
X1617 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1618 a_20863_n2724# vss a_20863_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1619 dac_3v_column_0[7].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[7].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1620 dvss a_n55547_n16609# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1621 dac_3v_column_odd_0[3].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_odd_0[3].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1622 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1623 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1624 dac_3v_column_odd_0[7].out1_0_0 dac_3v_8bit_0/b0b a_22563_n20019# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1625 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1626 dac_3v_column_0[1].out1_0_1 dac_3v_8bit_0/b0a a_25577_n6160# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1627 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1628 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1629 bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1630 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C a_n53615_n20961# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1631 vdd dac_3v_8bit_0/b6b dac_3v_8bit_0/b6a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1632 dac_3v_column_odd_0[0].out1_0_1 dac_3v_8bit_0/b0b a_25577_n5095# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1633 a_31412_n19346# dac_3v_8bit_0/b0a dac_3v_column_odd_0[7].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1634 a_23170_n15082# dac_3v_8bit_0/b1b dac_3v_column_odd_0[5].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1635 a_26891_n15082# dac_3v_8bit_0/b0a dac_3v_column_odd_0[5].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1636 bias_0.bi__pmirr_0.gate bias_0.bi__amplifier_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X1637 level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X1638 dac_3v_column_odd_0[1].out4 dac_3v_8bit_0/b4a dac_3v_column_odd_0[1].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1639 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1640 dac_3v_column_0[7].dum1_in dac_3v_column_0[7].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1641 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1642 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1643 a_22370_n12950# dac_3v_8bit_0/b0a dac_3v_column_odd_0[4].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1644 a_31605_n10424# dac_3v_column_odd_0[3].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1645 bandgap_0.bg__pnp_group_0.eg dvss a_n31275_n477# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1646 dvss level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1647 vdd a_14987_n11444# follower_amp_0.pdrv1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X1648 dvss a_n55047_n18669# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output6.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1649 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1650 a_29905_n17214# dac_3v_8bit_0/b0b dac_3v_column_odd_0[6].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1651 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1652 dac_3v_column_0[6].res1_in a_22370_n16147# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1653 a_20863_n10185# vdd a_20863_n10185# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1654 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1655 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1656 dac_3v_column_0[6].out1_0_2 dac_3v_8bit_0/b0a a_28591_n16820# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1657 a_20156_n2566# vdd a_20024_n2963# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1658 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1659 a_28398_n4422# a_29905_n4422# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1660 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1661 dac_3v_column_odd_0[1].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[1].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1662 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1663 a_28398_n10818# dac_3v_8bit_0/b0a dac_3v_column_odd_0[3].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1664 a_20156_n11094# vdd a_20156_n11094# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1665 a_23877_n10818# dac_3v_8bit_0/b0a dac_3v_column_odd_0[3].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1666 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1667 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1668 a_25384_n20410# a_26891_n20410# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1669 dvdd bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbp dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1670 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1671 follower_amp_0.ndrv a_13761_n11418# vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1672 vdd level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b7b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1673 testbuffer_0.tb__mux_0.tbm__passgate_0.en a_n54221_n16635# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1674 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1675 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1676 dac_3v_column_0[7].out_3 dac_3v_8bit_0/b3b dac_3v_column_0[7].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1677 a_27084_n21083# a_28591_n21083# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1678 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1679 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1680 a_28591_n12556# a_30098_n12556# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1681 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1682 dac_3v_column_0[7].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_0[7].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1683 dac_3v_column_0[4].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[4].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1684 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1685 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1686 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.X a_n55405_n20961# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1687 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1688 a_23170_n20686# vss a_22563_n21083# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1689 a_20156_n17490# vss dac_3v_column_odd_0[6].dum_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1690 testbuffer_0.tb__mux_0.tbm__passgate_5.en a_n53523_n22049# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1691 a_28398_n2290# vdd a_28398_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1692 a_26891_n11883# dac_3v_8bit_0/b0a dac_3v_column_0[4].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1693 vss follower_amp_0.nbias follower_amp_0.vcomn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1694 a_31412_n4422# dac_3v_column_odd_0[0].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1695 dac_3v_column_0[2].out1_0_0 dac_3v_8bit_0/b0b a_22563_n8292# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1696 a_26891_n20410# vdd a_26891_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1697 a_n23157_n925# a_n24701_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1698 a_29905_n16147# dac_3v_8bit_0/b0a dac_3v_column_0[6].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1699 dvss a_23802_3107# a_23802_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1700 a_22370_n20410# vss a_22370_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1701 dac_3v_column_odd_0[2].out_5 dac_3v_8bit_0/b5b dac_3v_column_odd_0[2].out4 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1702 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1703 dvss level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b6b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1704 a_33112_n21083# a_33112_n21083# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1705 dac_3v_column_odd_0[3].out4 dac_3v_8bit_0/b4a dac_3v_column_0[3].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1706 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1707 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1708 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1709 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1710 level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=2.1e+11p pd=2.06e+06u as=0p ps=0u w=750000u l=500000u
X1711 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1712 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1713 dvss a_22174_3107# a_22174_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1714 dvss dvss bandgap_0.bg__pnp_group_0.eg sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=1
X1715 vdd level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1716 a_22370_n4422# a_23877_n4422# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1717 a_28398_n14015# dac_3v_8bit_0/b0b dac_3v_column_0[5].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X1718 dvss a_27058_2206# level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X1719 level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1720 a_26891_n4422# dac_3v_8bit_0/b0b dac_3v_column_odd_0[0].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1721 dvss a_29626_3404# a_29264_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.2375e+12p ps=1.065e+07u w=1.5e+06u l=500000u
X1722 vdd dac_3v_8bit_0/b4a dac_3v_8bit_0/b4b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1723 a_31412_n2290# vdd a_31412_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1724 a_33719_n17490# vss a_33719_n17490# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1725 a_25577_n13623# a_27084_n13623# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1726 vdd dac_3v_8bit_0/b1a dac_3v_8bit_0/b1b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1727 a_22370_n14015# a_23877_n14015# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1728 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1729 dac_3v_column_0[6].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_0[6].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1730 a_20156_n16423# vdd dac_3v_column_0[6].dum1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1731 dac_3v_column_0[3].out1_0_3 dac_3v_8bit_0/b0b a_30098_n10424# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1732 dac_3v_column_0[3].out1_0_1 dac_3v_8bit_0/b0a a_24070_n10424# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1733 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1734 dvdd testbuffer_0.tb__mux_0.tbm__passgate_0.en a_n47185_n15278# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1735 a_34148_2837# a_34510_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X1736 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1737 dac_3v_column_0[6].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[6].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1738 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1739 dac_3v_column_odd_0[0].out0_2 dac_3v_8bit_0/b3a dac_3v_column_odd_0[0].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1740 a_34426_n18713# vss a_34426_n18713# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1741 dvdd a_n55547_n19873# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1742 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1743 dac_3v_8bit_0/b3a level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1744 dvss dac_3v_8bit_0/b0b dac_3v_8bit_0/b0a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1745 dvss dac_3v_8bit_0/b1a dac_3v_8bit_0/b1b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1746 dac_3v_column_0[7].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[7].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1747 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=1e+06u
X1748 testbuffer_0.tb__mux_0.tbm__passgate_6.en a_n54443_n22593# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1749 a_33719_n5763# vss a_33719_n5763# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1750 dac_3v_column_odd_0[2].out1_0_3 dac_3v_8bit_0/b0b a_31605_n9359# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1751 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1752 dac_3v_column_odd_0[7].dum_out1 vss a_34426_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1753 dvdd a_n53983_n17697# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1754 dvss a_34510_3404# a_34148_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1755 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1756 w_n19679_n3822# w_n19679_n3822# dvdd dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1757 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1758 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1759 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1760 a_23877_n5487# a_25384_n5487# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1761 vss a_13761_n11418# a_13761_n11418# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1762 dac_3v_column_odd_0[5].dum_in0 vdd a_34426_n15516# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1763 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n55353_n19355# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1764 dac_3v_column_0[4].dum1_in dac_3v_column_0[4].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1765 a_n32750_n1665# a_n31275_n2597# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1766 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1767 a_30098_n14688# a_31605_n14688# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1768 a_25384_n8686# a_26891_n8686# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1769 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1770 dac_3v_column_odd_0[5].out1_0_0 dac_3v_8bit_0/b0a a_22563_n15755# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1771 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inp bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1772 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1773 dac_3v_column_odd_0[5].out_3 dac_3v_8bit_0/b3a dac_3v_column_odd_0[5].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1774 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X a_n55547_n16609# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1775 vhigh dac_3v_8bit_0/b0a dac_3v_column_0[0].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1776 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1777 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1778 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1779 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1780 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1781 dac_3v_column_odd_0[1].dum_in0 vss a_34426_n6988# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1782 bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1783 dac_3v_column_odd_0[7].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_odd_0[7].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1784 a_23877_n11883# a_25384_n11883# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1785 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1786 a_23170_n15082# dac_3v_8bit_0/b1b dac_3v_column_odd_0[5].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1787 dac_3v_column_0[2].dum1_in dac_3v_column_0[2].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1788 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1789 dac_3v_8bit_0/b2a level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1790 a_n32750_n3785# a_n31275_n4717# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1791 a_31942_2371# a_31942_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1792 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1793 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1794 a_23877_n3355# dac_3v_8bit_0/b0a dac_3v_column_0[0].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X1795 a_23877_n14015# dac_3v_8bit_0/b0b dac_3v_column_0[5].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1796 testbuffer_0.tb__mux_0.tbm__passgate_6.en a_n54443_n22593# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1797 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1798 a_25384_n6554# dac_3v_8bit_0/b0b dac_3v_column_odd_0[1].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1799 a_n55547_n19873# in[1] dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1800 a_29905_n3355# a_31412_n3355# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1801 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X a_n55547_n16609# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1802 bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate a_n42353_11671# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X1803 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output4.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1804 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1805 vdd a_28686_2206# level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X1806 dac_3v_column_0[1].out1_0_3 dac_3v_8bit_0/b0b a_31605_n6160# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1807 dac_3v_column_odd_0[7].out1_0_2 dac_3v_8bit_0/b0a a_27084_n20019# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1808 dac_3v_column_0[1].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[1].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1809 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1810 a_n53645_n19873# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1811 dac_3v_column_odd_0[2].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_odd_0[2].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1812 dvdd bias_0.bi__pmirr_0.gate a_n40589_11447# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X1813 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbp dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1814 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1815 dac_3v_8bit_0/b5b dac_3v_8bit_0/b5a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1816 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1817 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1818 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n53983_n17697# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1819 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1820 dac_3v_column_0[5].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_0[5].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1821 dac_3v_column_odd_0[4].out1_0_1 dac_3v_8bit_0/b0b a_24070_n13623# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1822 dac_3v_column_odd_0[3].dum_out1 vdd a_34426_n12317# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1823 a_25577_n8292# a_27084_n8292# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1824 level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1825 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1826 dac_3v_column_0[6].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[6].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1827 dac_3v_column_odd_0[4].out_5 dac_3v_8bit_0/b5b dac_3v_column_odd_0[5].out4 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1828 a_23170_n10818# dac_3v_8bit_0/b1a dac_3v_column_odd_0[3].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1829 dac_3v_column_odd_0[2].res_in1 vdd a_20863_n9120# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1830 a_31412_n15082# dac_3v_column_odd_0[5].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1831 dac_3v_column_odd_0[4].res_in1 a_22370_n12950# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1832 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n54713_n20729# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1833 level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1834 a_26891_n12950# dac_3v_8bit_0/b0b dac_3v_column_odd_0[4].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1835 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1836 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1837 a_28398_n2724# vss a_28398_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1838 dac_3v_column_odd_0[0].out4 dac_3v_8bit_0/b4b dac_3v_column_odd_0[0].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1839 a_22370_n12950# dac_3v_8bit_0/b0b dac_3v_column_odd_0[4].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1840 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1841 dac_3v_column_odd_0[2].out_5 dac_3v_8bit_0/b6a dac_3v_column_odd_0[2].in_5 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1842 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbp dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1843 testbuffer_0.tb__mux_0.tbm__passgate_1.en a_n54221_n17179# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1844 dac_3v_column_0[5].out1_0_2 dac_3v_8bit_0/b0b a_27084_n14688# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1845 a_29905_n6554# dac_3v_8bit_0/b0a dac_3v_column_odd_0[1].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1846 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1847 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1848 a_23802_3107# b6 dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X1849 dvss level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1850 a_23170_n2566# vss a_23170_n2566# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1851 dac_3v_column_0[7].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_0[7].res1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X1852 a_33719_n4698# vdd dac_3v_column_odd_0[0].res_out1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X1853 follower_amp_0.vcomn2 dac_out a_16155_n11444# vss sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1854 dac_3v_column_0[4].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[4].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1855 dvss a_n21740_n3691# bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1856 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1857 a_28591_n20019# a_30098_n20019# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1858 a_31412_n20844# vss a_31412_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1859 dac_3v_column_odd_0[0].dum_in1 dac_3v_column_odd_0[0].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1860 a_n47950_6120# bias_0.bi__amplifier_0.bias dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1861 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1862 testbuffer_0.tb__mux_0.tbm__passgate_4.en a_n55233_n20443# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1863 dvss dac_3v_8bit_0/b5a dac_3v_8bit_0/b5b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1864 dac_3v_column_odd_0[0].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[0].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1865 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1866 a_21663_n20686# vss a_21663_n20686# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1867 dac_3v_column_0[3].out1_0_3 dac_3v_8bit_0/b0a a_30098_n10424# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1868 dac_3v_column_0[7].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[7].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1869 a_28398_n17214# a_29905_n17214# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1870 a_31412_n2724# vss a_31412_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1871 dac_3v_column_odd_0[0].out1_0_1 dac_3v_8bit_0/b0b a_24070_n5095# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1872 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1873 a_n53925_n19873# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n53645_n19873# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1874 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1875 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.X a_n55405_n20961# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1876 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1877 a_33719_n14291# vdd a_33719_n14291# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1878 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1879 dac_3v_column_0[0].out1_0_3 dac_3v_8bit_0/b0b a_30098_n4028# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1880 dac_3v_column_odd_0[0].out_5 dac_3v_8bit_0/b6a dac_3v_column_odd_0[2].in_5 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1881 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1882 a_27691_n20686# vss a_27084_n21083# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1883 dvdd a_n54221_n16635# testbuffer_0.tb__mux_0.tbm__passgate_0.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1884 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1885 a_33570_2206# a_33570_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X1886 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n47185_n24233# inp[7] dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1887 dac_3v_8bit_0/b2a level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1888 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1889 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output8.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1890 dac_3v_8bit_0/b2a level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1891 dac_3v_column_odd_0[4].dum_in0 vss a_34426_n13384# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1892 a_23802_2206# a_23802_2371# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X1893 a_20863_n3789# vdd a_20863_n3789# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1894 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1895 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1896 a_22370_n2724# vss a_22370_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1897 dac_3v_column_0[6].out1_0_0 dac_3v_8bit_0/b0b a_22563_n16820# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1898 a_20863_n14449# vdd a_20863_n14449# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1899 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1900 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1901 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1902 a_n55353_n19355# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1903 a_34426_n15516# vdd a_34426_n15516# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1904 dac_3v_column_odd_0[3].out1_0_1 dac_3v_8bit_0/b0a a_25577_n11491# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1905 dac_3v_column_0[0].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_0[0].res1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1906 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output6.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1907 dac_3v_column_0[2].res1_in vss a_20863_n8053# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=500000u
X1908 a_31412_n16147# dac_3v_8bit_0/b0a dac_3v_column_0[6].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1909 a_22370_n10818# a_23877_n10818# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1910 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1911 dvss a_26370_3404# a_26008_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.2375e+12p ps=1.065e+07u w=1.5e+06u l=500000u
X1912 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1913 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1914 dac_3v_column_odd_0[0].out1_0_2 dac_3v_8bit_0/b0a a_27084_n5095# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1915 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1916 a_23170_n19346# dac_3v_8bit_0/b1a dac_3v_column_odd_0[7].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1917 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1918 dac_3v_column_odd_0[5].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[5].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1919 a_34426_n6988# vss a_34426_n6988# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1920 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inn bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1921 dvss dac_3v_8bit_0/b2a dac_3v_8bit_0/b2b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1922 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1923 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1924 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1925 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1926 a_29905_n14015# dac_3v_8bit_0/b0b dac_3v_column_0[5].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1927 vdd level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1928 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1929 a_29264_2837# a_29626_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1930 dac_3v_column_odd_0[5].out1_0_1 dac_3v_8bit_0/b0b a_25577_n15755# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1931 dac_3v_column_odd_0[7].dum_in1 dac_3v_column_odd_0[7].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1932 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1933 dvdd a_28686_3107# a_29626_3404# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X1934 a_23877_n2290# a_25384_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1935 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1936 dvss level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b1a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1937 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1938 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/muxout dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X1939 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1940 a_30098_n11491# a_31605_n11491# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1941 dac_3v_column_odd_0[1].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_odd_0[1].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1942 bias_0.bi__amplifier_0.inn a_n20841_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1943 dvss a_25430_3107# a_26370_3404# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X1944 dac_3v_8bit_0/b7b level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1945 a_20156_n18555# vdd a_20156_n18555# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X1946 dac_3v_column_odd_0[5].out4 dac_3v_8bit_0/b4a dac_3v_column_0[5].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1947 a_20156_n7895# vdd a_20156_n7895# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1948 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1949 a_28398_n18279# dac_3v_8bit_0/b0a dac_3v_column_0[7].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1950 dac_3v_column_odd_0[6].dum_in1 dac_3v_column_odd_0[6].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1951 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1952 a_23877_n18279# dac_3v_8bit_0/b0a dac_3v_column_0[7].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X1953 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1954 dac_3v_column_odd_0[6].res_in1 a_22563_n17887# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1955 dvdd bias_0.bi__amplifier_0.mirr bias_0.bi__amplifier_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=6.32e+06u w=500000u l=1e+07u
X1956 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1957 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1958 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1959 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1960 sbamuxm4_0/vb[2] a_n32029_10936# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1961 dvss testbuffer_0.tb__mux_0.tbm__passgate_5.en a_n48623_n21248# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1962 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1963 dvdd a_n55547_n16609# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1964 dac_3v_column_0[5].out1_0_3 dac_3v_8bit_0/b0b a_30098_n14688# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1965 dac_3v_column_0[5].out1_0_1 dac_3v_8bit_0/b0a a_24070_n14688# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1966 dac_3v_column_0[4].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[4].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1967 dac_3v_column_0[2].out1_0_1 dac_3v_8bit_0/b0a a_24070_n8292# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X1968 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1969 dac_3v_column_odd_0[3].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_odd_0[3].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1970 dac_3v_column_odd_0[2].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[2].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X1971 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1972 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1973 dvss a_27058_3107# a_27058_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1974 a_20863_n11252# vss a_20863_n11252# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X1975 dac_3v_column_odd_0[1].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[1].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1976 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1977 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1978 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1979 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n54441_n21531# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1980 a_31412_n10818# dac_3v_8bit_0/b0b dac_3v_column_odd_0[3].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X1981 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1982 a_25384_n19346# dac_3v_8bit_0/b0a dac_3v_column_odd_0[7].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1983 dac_3v_column_odd_0[4].out_5 dac_3v_8bit_0/b6a dac_3v_column_odd_0[6].in_5 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1984 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1985 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1986 vdd level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b2a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1987 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1988 dac_3v_column_odd_0[7].res_in1 vss a_20863_n19780# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X1989 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1990 dvdd bias_0.bi__pmirr_0.gate a_n40589_12567# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X1991 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1992 testbuffer_0.tb__mux_0.tbm__passgate_1.en a_n54221_n17179# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1993 dvss a_34510_3404# a_34148_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1994 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1995 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1996 a_33719_n14291# vss a_33719_n14291# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X1997 a_25577_n10424# a_27084_n10424# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X1998 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1999 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2000 a_22752_2837# a_23114_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2001 a_28398_n9751# dac_3v_8bit_0/b0a dac_3v_column_0[3].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2002 a_26891_n9751# a_28398_n9751# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2003 sbamuxm4_0/vb[1] a_n32029_11780# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X2004 dvss testbuffer_0.tb__mux_0.tbm__passgate_7.en a_n48623_n24233# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X2005 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2006 dac_3v_column_odd_0[3].out0_2 dac_3v_8bit_0/b3b dac_3v_column_odd_0[3].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2007 dvss level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b0b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2008 dac_3v_column_odd_0[4].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[4].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2009 vdd level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b4a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2010 a_34426_n9120# vdd a_34426_n9120# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2011 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
D5 dvss b3 sky130_fd_pr__diode_pw2nd_05v5
X2012 dac_3v_column_odd_0[6].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[6].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2013 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2014 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2015 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2016 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2017 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2018 dvss a_23114_3404# a_22752_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2019 vdd dac_3v_8bit_0/b5a dac_3v_8bit_0/b5b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2020 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2021 dac_3v_column_odd_0[1].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_odd_0[1].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2022 a_n27017_n925# a_n27403_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X2023 vss follower_amp_0.nbias follower_amp_0.vcomn2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2024 dac_3v_column_odd_0[3].out4 dac_3v_8bit_0/b4a dac_3v_column_odd_0[3].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2025 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2026 dac_3v_column_0[1].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[1].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2027 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2028 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2029 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2030 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X2031 dvdd a_n54221_n17179# testbuffer_0.tb__mux_0.tbm__passgate_1.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2032 a_25384_n5487# a_26891_n5487# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2033 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2034 dac_3v_column_odd_0[5].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[5].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2035 a_22370_n6554# dac_3v_8bit_0/b0a dac_3v_column_odd_0[1].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2036 dac_3v_8bit_0/b7a dac_3v_8bit_0/b7b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2037 dac_3v_column_odd_0[1].res_in1 a_22370_n6554# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2038 dac_3v_column_0[4].out1_0_0 dac_3v_8bit_0/b0a a_22563_n12556# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2039 dac_3v_column_odd_0[2].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_odd_0[2].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2040 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2041 dac_3v_8bit_0/b6b level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2042 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2043 a_31412_n9751# dac_3v_8bit_0/b0a dac_3v_column_0[3].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2044 a_29905_n7619# a_31412_n7619# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2045 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2046 dac_3v_column_odd_0[7].res_in0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[7].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=500000u
X2047 dac_3v_column_0[4].out_3 dac_3v_8bit_0/b3a dac_3v_column_0[4].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2048 dac_3v_column_0[0].dum0_in vss a_34426_n3789# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2049 a_n54657_n18785# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n54937_n18785# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2050 dvss level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b1a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2051 dac_3v_column_0[6].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_0[6].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2052 dac_3v_column_odd_0[5].out1_0_3 dac_3v_8bit_0/b0b a_31605_n15755# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2053 dac_3v_column_odd_0[2].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[2].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2054 a_33719_n2566# vss vhigh vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2055 dac_3v_column_odd_0[3].out1_0_2 dac_3v_8bit_0/b0b a_28591_n11491# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2056 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2057 bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X2058 testbuffer_0.tb__mux_0.tbm__passgate_5.en a_n53523_n22049# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2059 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2060 a_n48347_n24233# a_n48623_n24233# dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X2061 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2062 sbamuxm4_0/vb[4] a_n32029_8404# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X2063 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2064 a_25430_2371# a_26008_2837# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.142e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=1e+06u
X2065 dac_3v_column_odd_0[7].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[7].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2066 bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__pmirr_0.vbn dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2067 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2068 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2069 a_25384_n3355# dac_3v_8bit_0/b0b dac_3v_column_0[0].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2070 dac_3v_column_odd_0[0].res_in1 vss a_20863_n4856# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2071 a_34426_n5921# vdd a_34426_n5921# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2072 a_27084_n7227# a_28591_n7227# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2073 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2074 a_n32750_1515# dvss bandgap_0.bg__pnp_group_0.eg dvss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X2075 dac_3v_column_0[6].out1_0_2 dac_3v_8bit_0/b0a a_27084_n16820# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2076 vdd dac_3v_8bit_0/b7b dac_3v_8bit_0/b7a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2077 dac_3v_8bit_0/b6b level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2078 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2079 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2080 sbamuxm4_0/ibp[0] bias_0.bi__pmirr_0.gate a_n42353_12119# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X2081 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2082 dac_3v_column_0[1].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_0[1].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2083 dvss dac_3v_8bit_0/b6b dac_3v_8bit_0/b6a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2084 a_23170_n6554# dac_3v_8bit_0/b1b dac_3v_column_odd_0[1].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2085 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2086 level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2087 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2088 dac_3v_column_0[3].out1_0_1 dac_3v_8bit_0/b0b a_24070_n10424# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2089 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2090 dac_3v_column_odd_0[2].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[2].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2091 dvss in[2] a_n55681_n22593# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X2092 dvss level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b5a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2093 dac_3v_column_0[1].res1_in vdd a_20863_n5921# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2094 follower_amp_0.vcomn1 dac_3v_8bit_0/out_unbuf follower_amp_0.pdrv1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2095 dac_3v_column_0[7].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_0[7].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2096 dac_3v_column_0[4].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[4].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2097 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2098 bandgap_0.bg__pnp_group_0.eg dvss a_n31275_n2597# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2099 dac_3v_column_0[1].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_0[1].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2100 dac_3v_column_0[5].out1_0_3 dac_3v_8bit_0/b0a a_30098_n14688# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2101 a_31412_n11883# dac_3v_column_odd_0[3].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2102 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2103 a_26008_2837# a_26370_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2104 dac_3v_column_0[7].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[7].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2105 dac_3v_column_odd_0[0].out_3 dac_3v_8bit_0/b3a dac_3v_column_odd_0[0].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2106 dvdd a_25430_3107# a_26370_3404# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X2107 a_30098_n5095# a_31605_n5095# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2108 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2109 sbamuxm4_0/vb[3] a_n32029_9248# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X2110 dac_3v_column_odd_0[0].out_5 dac_3v_8bit_0/b5b dac_3v_column_odd_0[1].out4 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2111 a_22563_n18952# a_24070_n18952# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2112 a_28398_n20410# vss a_28398_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2113 a_29905_n3355# dac_3v_8bit_0/b0a dac_3v_column_0[0].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2114 a_23170_n8686# dac_3v_8bit_0/b1b dac_3v_column_odd_0[2].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2115 dac_3v_8bit_0/b2a level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2116 dac_3v_column_0[0].out1_0_2 dac_3v_8bit_0/b0a a_28591_n4028# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2117 a_20156_n4698# vdd a_20156_n4698# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2118 a_28398_n15082# dac_3v_8bit_0/b0a dac_3v_column_odd_0[5].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2119 a_20156_n15358# vdd a_20156_n15358# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2120 a_28398_n7619# dac_3v_8bit_0/b0b dac_3v_column_0[2].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2121 a_24677_n2566# vss a_24677_n2566# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2122 a_29198_n2566# vss a_28591_n2963# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2123 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2124 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._17_.X a_n53523_n22049# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2125 a_23877_n15082# dac_3v_8bit_0/b0a dac_3v_column_odd_0[5].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2126 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2127 bandgap_0.bg__pnp_group_0.eg dvss a_n31275_n4717# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2128 level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2129 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2130 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2131 dvss a_n54221_n16635# testbuffer_0.tb__mux_0.tbm__passgate_0.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2132 a_30892_2837# a_30314_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=1e+06u
X2133 dac_3v_column_odd_0[4].out1_0_3 dac_3v_8bit_0/b0a a_31605_n13623# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2134 a_20156_n11094# vss dac_3v_column_odd_0[3].dum_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2135 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2136 dac_3v_column_odd_0[7].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_odd_0[7].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2137 a_28398_n14015# a_29905_n14015# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2138 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2139 a_22174_2206# a_22174_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X2140 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2141 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2142 dac_3v_column_odd_0[0].out1_0_1 dac_3v_8bit_0/b0a a_25577_n5095# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2143 a_20156_n19622# vss a_20156_n19622# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2144 dvdd in[2] a_n55681_n22593# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X2145 dac_3v_column_odd_0[2].out4 dac_3v_8bit_0/b4b dac_3v_column_0[2].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2146 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2147 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2148 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2149 dac_3v_column_0[0].out1_0_3 dac_3v_8bit_0/b0a a_31605_n4028# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2150 dac_3v_column_odd_0[2].res_out1 dac_3v_column_odd_0[2].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2151 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2152 dac_3v_column_0[3].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[3].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2153 a_31412_n7619# dac_3v_8bit_0/b0b dac_3v_column_0[2].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2154 a_n41084_8994# bias_0.bi__nmirr_0.gate_n dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X2155 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X a_n55547_n16609# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2156 dvss dac_3v_8bit_0/b0b dac_3v_8bit_0/b0a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2157 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X2158 dvdd bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2159 dac_3v_column_odd_0[1].out1_0_3 dac_3v_8bit_0/b0a a_30098_n7227# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2160 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2161 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2162 vdd dac_3v_8bit_0/b0b dac_3v_8bit_0/b0a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2163 dac_3v_column_odd_0[7].out1_0_2 dac_3v_8bit_0/b0b a_27084_n20019# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2164 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n55547_n19873# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2165 a_24070_n21083# a_25577_n21083# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2166 a_34426_n12317# vdd a_34426_n12317# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2167 dac_3v_column_0[7].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[7].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2168 dac_3v_column_0[2].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[2].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2169 a_27058_2371# a_27058_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2170 a_20156_n12159# vdd a_20156_n12159# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2171 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2172 dac_3v_column_0[0].out1_0_0 dac_3v_8bit_0/b0a a_22563_n4028# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2173 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2174 dac_3v_column_odd_0[5].out1_0_2 dac_3v_8bit_0/b0a a_28591_n15755# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2175 a_28398_n11883# dac_3v_8bit_0/b0a dac_3v_column_0[4].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2176 dac_3v_column_odd_0[1].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[1].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2177 dvss a_30314_2206# level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X2178 a_23877_n11883# dac_3v_8bit_0/b0a dac_3v_column_0[4].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2179 a_22370_n7619# dac_3v_8bit_0/b0b dac_3v_column_0[2].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2180 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2181 level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X2182 dac_3v_column_0[6].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[6].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2183 a_25384_n15082# a_26891_n15082# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2184 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2185 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2186 a_23877_n20410# vdd a_23877_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2187 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2188 vdd level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2189 a_20156_n8962# vss dac_3v_column_odd_0[2].dum_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2190 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2191 a_27084_n15755# a_28591_n15755# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2192 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2193 dvss a_n54221_n17179# testbuffer_0.tb__mux_0.tbm__passgate_1.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2194 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2195 dac_3v_column_0[7].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_0[7].res1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X2196 dac_3v_column_0[4].out1_0_1 dac_3v_8bit_0/b0b a_25577_n12556# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2197 dac_3v_8bit_0/b7a dac_3v_8bit_0/b7b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2198 dac_3v_8bit_0/b3a level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2199 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2200 dac_3v_column_odd_0[6].out_3 dac_3v_8bit_0/b3b dac_3v_column_odd_0[6].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2201 a_33570_3107# b0 dvss dvss sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X2202 a_25384_n20844# vss a_25384_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2203 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2204 dac_3v_column_odd_0[6].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[6].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2205 a_n32750_1515# a_n31275_583# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X2206 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2207 a_25384_n2290# a_26891_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2208 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2209 a_21663_n20686# vdd a_21663_n20686# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2210 dac_3v_column_odd_0[4].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_odd_0[4].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2211 a_20863_n19780# vdd a_20863_n19780# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2212 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X2213 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2214 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2215 dac_3v_8bit_0/b5b dac_3v_8bit_0/b5a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2216 dvss level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b0b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2217 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2218 dac_3v_column_odd_0[5].res_out1 dac_3v_column_odd_0[5].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2219 dac_3v_column_0[5].dum1_in dac_3v_column_0[5].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2220 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2221 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2222 dvss a_n53615_n20961# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2223 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2224 a_23170_n17214# dac_3v_8bit_0/b1b dac_3v_column_odd_0[6].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2225 dac_3v_column_odd_0[1].out1_0_1 dac_3v_8bit_0/b0b a_25577_n7227# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2226 dvss a_n55547_n16609# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2227 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2228 a_26891_n17214# dac_3v_8bit_0/b0a dac_3v_column_odd_0[6].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2229 dac_3v_column_0[5].res1_in a_22563_n14688# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2230 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbp dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2231 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2232 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n55681_n18241# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2233 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2234 a_27691_n20686# vdd a_27084_n21083# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2235 dvss a_33570_3107# a_33570_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2236 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2237 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2238 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2239 dvdd a_n54587_n22049# a_n54487_n21933# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2240 a_28398_n12950# dac_3v_8bit_0/b0b dac_3v_column_odd_0[4].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2241 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2242 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2243 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2244 a_20156_n5763# vss dac_3v_column_0[1].dum1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2245 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2246 a_33719_n18555# vdd dac_3v_column_odd_0[7].res_in0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2247 dac_3v_8bit_0/b2a level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2248 a_28398_n6554# a_29905_n6554# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2249 dac_3v_column_odd_0[5].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_odd_0[5].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2250 a_20156_n15358# vdd dac_3v_column_odd_0[5].dum_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2251 vss follower_amp_0.nbias follower_amp_0.nbias vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2252 dvss bias_0.bi__amplifier_0.bias a_n47950_6120# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X2253 vdd a_31942_2206# level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X2254 a_34426_n17648# vss a_34426_n17648# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2255 a_25384_n16147# dac_3v_8bit_0/b0a dac_3v_column_0[6].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2256 dac_3v_column_odd_0[5].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[5].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2257 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2258 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/muxout dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.48e+12p ps=2.574e+07u w=4e+06u l=4e+06u
X2259 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2260 dac_3v_column_0[6].res1_in vss a_20863_n16581# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2261 a_n25473_n925# a_n24315_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X2262 dvss a_23114_3404# a_22752_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2263 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2264 a_31412_n18279# dac_3v_8bit_0/b0b dac_3v_column_0[7].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2265 dac_3v_column_odd_0[7].out4 dac_3v_8bit_0/b4b dac_3v_column_odd_0[7].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2266 a_33719_n20686# vdd a_33719_n20686# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2267 dvss level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2268 a_22370_n19346# a_23877_n19346# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2269 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2270 bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2271 a_n55047_n18669# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2272 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2273 dvss level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2274 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2275 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2276 a_23170_n15082# dac_3v_8bit_0/b1a dac_3v_column_odd_0[5].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2277 vdd level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b6b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2278 a_n41084_9346# bias_0.bi__nmirr_0.gate_n dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X2279 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n53615_n20961# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2280 a_24380_2837# a_24742_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2281 a_20863_n20844# vdd a_20863_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2282 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2283 dac_3v_8bit_0/b6a dac_3v_8bit_0/b6b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2284 dac_3v_column_0[3].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[3].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2285 bias_0.bi__amplifier_0.bias bias_basis_current_0.bb__pmirr_0.vbp dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2286 a_28398_n4422# dac_3v_8bit_0/b0b dac_3v_column_odd_0[0].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2287 follower_amp_0.pdrv2 a_16155_n11444# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X2288 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2289 dac_3v_column_0[7].out0_2 dac_3v_8bit_0/b3b dac_3v_column_0[7].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2290 dac_3v_column_odd_0[1].res_in0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[1].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2291 a_32919_n2290# vss a_32919_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2292 a_31412_n6554# dac_3v_column_odd_0[1].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2293 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2294 dac_3v_column_odd_0[7].out1_0_3 dac_3v_8bit_0/b0b a_30098_n20019# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2295 a_n23132_n3629# bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvdd dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2296 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2297 level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X2298 dvss level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2299 dac_3v_column_odd_0[7].out1_0_1 dac_3v_8bit_0/b0a a_24070_n20019# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2300 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2301 dac_3v_column_0[0].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_0[0].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2302 dac_3v_column_0[7].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[7].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2303 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2304 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2305 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2306 dvss a_24742_3404# a_24380_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2307 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2308 a_33719_n6830# vdd a_33719_n6830# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2309 a_22370_n3355# dac_3v_8bit_0/b0a dac_3v_column_0[0].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2310 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2311 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2312 bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas bias_0.bi__nmirr_0.gate_n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2313 dac_3v_column_0[0].res1_in a_22370_n3355# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2314 a_28398_n10818# a_29905_n10818# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2315 dvss bias_0.bi__nmirr_0.gate_n dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2316 a_29905_n20410# vdd a_29905_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2317 dac_3v_column_odd_0[5].res_out1 dac_3v_8bit_0/b0a dac_3v_column_0[6].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2318 a_23877_n6554# dac_3v_8bit_0/b0b dac_3v_column_odd_0[1].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2319 a_23877_n2290# vss a_23877_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2320 a_22370_n6554# a_23877_n6554# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2321 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2322 a_23877_n12950# dac_3v_8bit_0/b0b dac_3v_column_odd_0[4].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2323 dac_3v_column_odd_0[2].out_3 dac_3v_8bit_0/b3b dac_3v_column_odd_0[2].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2324 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output7.A a_n55313_n22049# dvss dvss sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2325 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output6.A a_n54301_n18241# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2326 a_n48347_n15278# a_n48623_n15278# dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X2327 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2328 a_31412_n4422# dac_3v_8bit_0/b0b dac_3v_column_odd_0[0].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2329 dac_3v_column_0[1].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[1].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2330 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2331 a_22370_n16147# a_23877_n16147# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2332 dac_3v_column_0[5].out1_0_1 dac_3v_8bit_0/b0b a_24070_n14688# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2333 dac_3v_column_0[4].out1_0_3 dac_3v_8bit_0/b0b a_31605_n12556# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2334 a_23170_n6554# dac_3v_8bit_0/b2b dac_3v_column_odd_0[1].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2335 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2336 dac_3v_8bit_0/b2b dac_3v_8bit_0/b2a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2337 dac_3v_column_odd_0[0].out1_0_3 dac_3v_8bit_0/b0b a_31605_n5095# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2338 dac_3v_column_odd_0[2].out1_0_2 dac_3v_8bit_0/b0b a_27084_n9359# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2339 vdd dac_3v_8bit_0/b0b dac_3v_8bit_0/b0a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2340 dac_3v_column_0[4].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[4].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2341 a_32919_n20844# vdd a_32919_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2342 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2343 a_n40589_12343# bias_0.bi__pmirr_0.gate sbamuxm4_0/ibp[2] dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X2344 a_29264_2837# a_28686_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=1e+06u
X2345 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2346 a_26891_n18279# a_28398_n18279# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2347 dac_3v_column_0[6].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[6].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2348 a_33719_n7895# vss a_33719_n7895# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2349 dac_3v_column_odd_0[4].out_5 dac_3v_8bit_0/b6b dac_3v_column_odd_0[6].in_5 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2350 a_25384_n10818# dac_3v_8bit_0/b0b dac_3v_column_odd_0[3].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2351 a_27084_n4028# a_28591_n4028# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2352 testbuffer_0.tb__mux_0.tbm__passgate_7.en a_n53197_n22593# dvss dvss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X2353 a_22370_n4422# dac_3v_8bit_0/b0b dac_3v_column_odd_0[0].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2354 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2355 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2356 sbamuxm4_0/ibp[0] bias_0.bi__pmirr_0.gate a_n42353_11895# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X2357 sbamuxm4_0/ibn[0] bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[0] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2358 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2359 testbuffer_0.tb__mux_0.tbm__passgate_6.en a_n54443_n22593# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2360 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2361 a_25430_2371# a_25430_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2362 dac_3v_column_odd_0[6].dum_in0 vdd a_34426_n17648# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2363 dvdd a_n55547_n19873# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2364 dac_3v_column_0[0].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[0].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2365 a_30098_n16820# a_31605_n16820# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2366 level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2367 a_30705_n20686# vdd a_30098_n21083# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2368 a_24677_n20686# vss a_24070_n21083# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2369 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output5.A a_n54035_n19757# a_n53925_n19873# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2370 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2371 dvss level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b6b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2372 dac_3v_column_0[1].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[1].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2373 dac_3v_column_odd_0[6].res_out1 dac_3v_column_odd_0[6].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2374 dac_3v_column_odd_0[6].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[6].res_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2375 dac_3v_column_odd_0[1].out0_2 dac_3v_8bit_0/b3b dac_3v_column_odd_0[1].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2376 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2377 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2378 dac_3v_column_odd_0[3].out0_2 dac_3v_8bit_0/b3a dac_3v_column_odd_0[3].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2379 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2380 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2381 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2382 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 sbamuxm4_0/ibp[0] sbamuxm4_0/ibp[0] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=4e+06u
X2383 dac_3v_column_0[1].out_3 dac_3v_8bit_0/b3b dac_3v_column_0[1].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2384 bias_0.bi__pmirr_0.gate bias_0.bi__amplifier_0.inn bias_0.bi__amplifier_0.diff dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X2385 vdd level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2386 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2387 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2388 a_33719_n18555# vss dac_3v_column_odd_0[7].res_in0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2389 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2390 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2391 vhigh dac_3v_column_0[0].dum0_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2392 a_23170_n17214# dac_3v_8bit_0/b1b dac_3v_column_odd_0[6].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2393 dac_3v_column_0[3].dum1_in dac_3v_column_0[3].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2394 a_n53553_n18785# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2395 level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2396 dac_3v_column_0[1].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[1].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2397 dac_3v_column_0[1].out1_0_2 dac_3v_8bit_0/b0b a_27084_n6160# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2398 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2399 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2400 dvss a_n54945_n17689# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.X dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2401 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2402 dac_3v_column_odd_0[3].dum_in1 dac_3v_column_odd_0[3].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2403 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2404 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2405 a_33719_n20686# vss a_33719_n20686# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2406 a_30705_n2566# vdd a_30098_n2963# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2407 a_33719_n13226# vdd a_33719_n13226# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2408 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2409 dvss dac_3v_8bit_0/b1a dac_3v_8bit_0/b1b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2410 bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas bias_0.bi__nmirr_0.gate_n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2411 dvdd a_n53197_n19329# testbuffer_0.tb__mux_0.tbm__passgate_2.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2412 dac_3v_column_odd_0[3].res_in1 a_22563_n11491# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2413 a_n25087_n925# a_n26245_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X2414 testbuffer_0.tb__mux_0.tbm__passgate_7.en a_n53197_n22593# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2415 dvss level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b7b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2416 dac_3v_column_0[2].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[2].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2417 dac_3v_8bit_0/b4b dac_3v_8bit_0/b4a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2418 dac_3v_column_0[3].out1_0_3 dac_3v_8bit_0/b0a a_31605_n10424# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2419 testbuffer_0.tb__mux_0.tbm__passgate_6.en a_n54443_n22593# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2420 a_20863_n2724# vdd a_20863_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2421 dvss bias_0.bi__pmirr_0.gate_cas dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2422 dac_3v_column_0[6].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_0[6].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2423 dac_3v_column_odd_0[5].out1_0_0 dac_3v_8bit_0/b0b a_22563_n15755# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2424 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2425 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2426 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.X a_n54443_n22593# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2427 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2428 a_33570_2206# a_33570_2371# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X2429 dac_3v_column_odd_0[3].res_in1 vdd a_20863_n11252# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X2430 bias_0.bi__pmirr_0.gate bias_0.bi__amplifier_0.inn bias_0.bi__amplifier_0.diff dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X2431 a_20156_n16423# vss a_20156_n16423# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2432 a_21663_n2566# vdd a_20863_n2290# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2433 dac_3v_column_odd_0[7].out1_0_3 dac_3v_8bit_0/b0a a_30098_n20019# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2434 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2435 dvss a_n55233_n20443# testbuffer_0.tb__mux_0.tbm__passgate_4.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2436 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2437 dac_3v_column_odd_0[1].res_in0 dac_3v_column_odd_0[1].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2438 a_34426_n8053# vss a_34426_n8053# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2439 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2440 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2441 vdd dac_3v_8bit_0/b2a dac_3v_8bit_0/b2b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2442 dac_3v_column_odd_0[1].out4 dac_3v_8bit_0/b4b dac_3v_column_odd_0[1].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2443 dvss a_30314_3107# a_30314_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2444 dac_3v_column_0[3].out0_1_1 dac_3v_8bit_0/b2a dac_3v_column_0[3].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2445 a_n54713_n20729# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2446 a_n53615_n20961# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2447 dac_3v_column_0[6].out1_0_2 dac_3v_8bit_0/b0b a_27084_n16820# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2448 dac_3v_8bit_0/b0b level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2449 a_31412_n15082# dac_3v_8bit_0/b0b dac_3v_column_odd_0[5].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2450 dac_3v_8bit_0/b4a level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2451 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2452 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2453 dvss level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2454 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2455 a_33719_n6830# vdd dac_3v_column_odd_0[1].res_out1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2456 sbamuxm4_0/ibn[1] bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[1] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2457 dac_3v_8bit_0/b6b level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2458 a_29905_n12950# dac_3v_8bit_0/b0b dac_3v_column_odd_0[4].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2459 a_n53825_n18785# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n53553_n18785# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2460 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2461 dac_3v_column_0[4].out1_0_2 dac_3v_8bit_0/b0a a_28591_n12556# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2462 dac_3v_column_0[2].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_0[2].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2463 dac_3v_column_odd_0[1].dum_in1 dac_3v_column_odd_0[1].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2464 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2465 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2466 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2467 dac_3v_column_odd_0[1].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[1].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2468 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2469 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2470 a_25384_n11883# a_26891_n11883# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2471 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2472 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2473 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2474 dac_3v_column_odd_0[5].out0_2 dac_3v_8bit_0/b3b dac_3v_column_odd_0[5].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2475 dac_3v_column_odd_0[3].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[3].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2476 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2477 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2478 a_27084_n12556# a_28591_n12556# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2479 dac_3v_column_odd_0[1].out1_0_1 dac_3v_8bit_0/b0b a_24070_n7227# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2480 dac_3v_column_odd_0[2].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[2].res_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2481 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.X a_n54443_n22593# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2482 dac_3v_column_odd_0[3].res_in0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[3].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2483 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2484 a_n46909_n18263# a_n47185_n18263# dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X2485 vdd level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
D6 dvss b1 sky130_fd_pr__diode_pw2nd_05v5
X2486 dvss dvss dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X2487 a_22370_n19346# dac_3v_8bit_0/b0a dac_3v_column_odd_0[7].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2488 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inp bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2489 a_n54345_n20265# a_n54072_n20437# a_n54114_n20411# dvss sky130_fd_pr__nfet_01v8 ad=1.07825e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2490 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output8.A a_n54441_n21531# a_n54691_n21255# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2491 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2492 a_29905_n20410# a_31412_n20410# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2493 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2494 dvss level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b7b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2495 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2496 dvdd a_n54221_n16635# testbuffer_0.tb__mux_0.tbm__passgate_0.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2497 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2498 dac_3v_column_0[3].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_0[3].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2499 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2500 a_31605_n21083# a_33112_n21083# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2501 a_20863_n16581# vdd a_20863_n16581# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2502 dac_3v_column_0[2].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[2].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2503 dvdd testbuffer_0.tb__mux_0.tbm__passgate_7.en a_n48623_n24233# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X2504 a_30705_n20686# vss a_30098_n21083# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2505 dac_3v_column_odd_0[4].res_in0 dac_3v_column_odd_0[4].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2506 dac_3v_column_odd_0[4].out1_0_1 dac_3v_8bit_0/b0a a_25577_n13623# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2507 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2508 dac_3v_column_0[5].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[5].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2509 a_31412_n11883# dac_3v_8bit_0/b0b dac_3v_column_0[4].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2510 dac_3v_column_odd_0[3].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_odd_0[3].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2511 bandgap_0.bg__pnp_group_0.eg dvss a_n31275_1643# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2512 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2513 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2514 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2515 a_22370_n12950# a_23877_n12950# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2516 a_23170_n10818# dac_3v_8bit_0/b2a dac_3v_column_odd_0[3].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2517 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2518 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2519 a_26891_n14015# dac_3v_8bit_0/b0a dac_3v_column_0[5].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2520 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2521 dac_3v_8bit_0/b6a dac_3v_8bit_0/b6b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2522 dac_3v_8bit_0/b0b level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2523 dac_3v_column_odd_0[1].out1_0_2 dac_3v_8bit_0/b0a a_27084_n7227# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2524 a_n21613_n925# a_n22771_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X2525 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n55353_n19355# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2526 a_n54035_n19757# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvss dvss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2527 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2528 a_22174_3107# b7 dvss dvss sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X2529 dac_3v_8bit_0/b2b dac_3v_8bit_0/b2a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2530 dac_3v_column_odd_0[6].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[6].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2531 dac_3v_8bit_0/b6a dac_3v_8bit_0/b6b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2532 a_33719_n4698# vss a_33719_n4698# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2533 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2534 dvss dac_3v_8bit_0/b4a dac_3v_8bit_0/b4b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2535 a_28591_n18952# a_30098_n18952# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2536 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2537 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2538 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2539 dac_3v_column_0[5].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[5].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2540 dac_3v_column_0[4].out0_2 dac_3v_8bit_0/b3b dac_3v_column_0[4].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2541 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2542 vdd dac_3v_8bit_0/b2a dac_3v_8bit_0/b2b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2543 dac_3v_column_0[1].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_0[1].res1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2544 a_33719_n13226# vss a_33719_n13226# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2545 a_28398_n8686# dac_3v_8bit_0/b0a dac_3v_column_odd_0[2].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2546 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2547 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2548 dvss a_27998_3404# a_27636_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2549 dac_3v_8bit_0/b0a dac_3v_8bit_0/b0b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2550 a_28398_n3355# a_29905_n3355# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2551 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2552 dac_3v_column_0[4].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_0[4].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2553 a_20156_n12159# vdd dac_3v_column_0[4].dum1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2554 a_26891_n8686# a_28398_n8686# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2555 vdd level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2556 dac_3v_column_0[4].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[4].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2557 dvss bias_0.bi__amplifier_0.bias bias_0.bi__amplifier_0.bias dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X2558 a_30098_n13623# a_31605_n13623# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2559 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2560 dvss a_22174_3107# a_22174_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2561 a_32520_2837# a_32882_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2562 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2563 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2564 dvss dac_3v_8bit_0/b1a dac_3v_8bit_0/b1b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2565 dac_3v_column_odd_0[6].out4 dac_3v_8bit_0/b4a dac_3v_column_0[6].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2566 vdd a_33570_2206# level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X2567 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2568 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2569 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n46909_n15278# inp[0] dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2570 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2571 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2572 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2573 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2574 level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2575 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n55547_n19873# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2576 dvss a_24742_3404# a_24380_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2577 dvss a_23802_2206# level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X2578 dvss level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2579 a_n54587_n22049# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2580 dac_3v_8bit_0/b3b dac_3v_8bit_0/b3a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2581 dac_3v_column_0[2].res1_in a_22370_n7619# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2582 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2583 dvss a_32882_3404# a_32520_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2584 dac_3v_column_odd_0[0].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[0].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2585 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2586 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n53983_n17697# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2587 a_26891_n6554# dac_3v_8bit_0/b0a dac_3v_column_odd_0[1].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2588 a_n54713_n20729# a_n54440_n20729# a_n54482_n20601# dvss sky130_fd_pr__nfet_01v8 ad=1.07825e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X2589 vhigh dac_3v_8bit_0/b0b dac_3v_column_0[0].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2590 a_31412_n8686# dac_3v_8bit_0/b0a dac_3v_column_odd_0[2].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2591 a_31412_n3355# vhigh vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2592 dac_3v_column_0[6].out1_0_3 dac_3v_8bit_0/b0b a_30098_n16820# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2593 dvdd a_n55353_n19355# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2594 dac_3v_column_0[6].out1_0_1 dac_3v_8bit_0/b0a a_24070_n16820# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2595 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2596 a_32919_n2290# vss a_34426_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2597 dac_3v_column_odd_0[4].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_odd_0[4].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2598 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2599 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2600 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._19_.A a_n53289_n21505# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2601 a_20863_n13384# vss a_20863_n13384# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2602 a_33719_n3631# vdd a_33719_n3631# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2603 dac_3v_column_odd_0[5].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_odd_0[5].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2604 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2605 dvdd a_n55547_n16609# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2606 dac_3v_column_odd_0[0].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[0].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2607 bias_0.bi__nmirr_0.gate_n bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2608 a_27084_n8292# a_28591_n8292# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2609 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbn dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2610 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2611 a_23877_n3355# dac_3v_8bit_0/b0b dac_3v_column_0[0].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2612 dac_3v_column_0[0].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_0[0].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2613 a_22370_n3355# a_23877_n3355# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2614 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2615 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2616 dac_3v_8bit_0/b1b dac_3v_8bit_0/b1a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2617 a_25384_n2290# vss a_25384_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2618 a_34426_n4856# vdd a_34426_n4856# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2619 dac_3v_column_0[7].dum1_in dac_3v_column_0[7].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2620 bandgap_0.bg__pnp_group_0.eg dvss a_n31275_n1537# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2621 dac_3v_column_0[0].out0_1_1 dac_3v_8bit_0/b2b dac_3v_column_0[0].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2622 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2623 dac_3v_column_odd_0[5].out1_0_2 dac_3v_8bit_0/b0a a_27084_n15755# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2624 dac_3v_column_odd_0[2].res_out1 dac_3v_8bit_0/b0a dac_3v_column_0[3].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=500000u
X2625 a_23170_n6554# dac_3v_8bit_0/b1a dac_3v_column_odd_0[1].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2626 dac_3v_8bit_0/b1b dac_3v_8bit_0/b1a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2627 a_n32750_2575# dvss bandgap_0.bg__pnp_group_0.eg dvss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X2628 vdd level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b6b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2629 dac_3v_column_odd_0[0].res_in1 a_22563_n5095# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2630 dvss a_25430_3107# a_25430_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2631 dac_3v_column_odd_0[0].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_odd_0[0].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2632 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2633 dac_3v_column_odd_0[6].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_odd_0[6].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2634 a_25384_n18279# dac_3v_8bit_0/b0b dac_3v_column_0[7].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2635 dac_3v_column_0[0].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_0[0].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2636 dac_3v_column_odd_0[3].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_odd_0[3].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2637 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2638 a_30314_2371# a_30314_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2639 dac_3v_column_odd_0[4].dum_out1 vdd a_34426_n14449# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2640 dac_3v_column_odd_0[4].out4 dac_3v_8bit_0/b4a dac_3v_column_odd_0[4].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2641 bandgap_0.bg__pnp_group_0.eg dvss a_n31275_n3657# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X2642 a_23877_n9751# dac_3v_8bit_0/b0a dac_3v_column_0[3].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2643 a_22563_n17887# a_24070_n17887# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2644 a_27084_n20019# a_28591_n20019# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2645 dvdd bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2646 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbn dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2647 dac_3v_column_odd_0[6].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[6].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2648 a_29905_n2290# vss a_29905_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2649 a_29198_n2566# vdd a_28591_n2963# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2650 dac_3v_column_0[0].out0_2 dac_3v_8bit_0/b3b dac_3v_column_0[0].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2651 a_29905_n9751# a_31412_n9751# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2652 dac_3v_8bit_0/b4a level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2653 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2654 a_n23543_n925# a_n22385_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X2655 follower_amp_0.pdrv1 a_14987_n11444# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2656 dvdd a_n54221_n17179# testbuffer_0.tb__mux_0.tbm__passgate_1.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2657 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2658 dac_3v_column_0[7].out0_2 dac_3v_8bit_0/b3a dac_3v_column_0[7].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2659 dac_3v_column_0[5].out1_0_3 dac_3v_8bit_0/b0a a_31605_n14688# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2660 a_26891_n17214# a_28398_n17214# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2661 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2662 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2663 dac_3v_column_odd_0[3].out_3 dac_3v_8bit_0/b3b dac_3v_column_odd_0[3].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2664 dac_3v_column_odd_0[7].out1_0_1 dac_3v_8bit_0/b0b a_24070_n20019# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2665 dac_3v_column_odd_0[4].out1_0_2 dac_3v_8bit_0/b0b a_28591_n13623# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2666 vlow dac_3v_column_odd_0[7].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2667 dac_3v_column_odd_0[3].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[3].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2668 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2669 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2670 dac_3v_column_0[5].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[5].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2671 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2672 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2673 vdd level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2674 dac_3v_8bit_0/b6a dac_3v_8bit_0/b6b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2675 dac_3v_8bit_0/b4a level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2676 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2677 a_24070_n9359# a_25577_n9359# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2678 dvdd a_n55233_n20443# testbuffer_0.tb__mux_0.tbm__passgate_4.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2679 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2680 a_26891_n19346# dac_3v_8bit_0/b0b dac_3v_column_odd_0[7].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2681 level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2682 a_20863_n9120# vss a_20863_n9120# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2683 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2684 dvss level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2685 a_22370_n19346# dac_3v_8bit_0/b0b dac_3v_column_odd_0[7].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2686 bias_0.bi__nmirr_0.gate_n bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X2687 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2688 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2689 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2690 dac_3v_column_odd_0[6].res_in0 dac_3v_column_odd_0[6].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2691 dac_3v_column_0[2].out1_0_3 dac_3v_8bit_0/b0a a_30098_n8292# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2692 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2693 a_32212_n2566# vdd a_31605_n2963# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2694 a_23170_n8686# dac_3v_8bit_0/b1a dac_3v_column_odd_0[2].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2695 a_28398_n19346# a_29905_n19346# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2696 vdd level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b5a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2697 dac_3v_8bit_0/b4a level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2698 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbp dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2699 a_24070_n15755# a_25577_n15755# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2700 dac_3v_column_0[2].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_0[2].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2701 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2702 dac_3v_column_0[4].out1_0_0 dac_3v_8bit_0/b0b a_22563_n12556# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2703 dac_3v_column_0[2].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_0[2].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2704 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2705 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2706 sbamuxm4_0/vb[2] a_n32029_10092# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X2707 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2708 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output5.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2709 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output8.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2710 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2711 dac_3v_column_odd_0[6].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[6].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2712 dac_3v_column_0[2].res1_in vdd a_20863_n8053# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2713 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 sbamuxm4_0/ibp[0] sbamuxm4_0/ibp[0] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2714 dac_3v_column_0[6].out1_0_3 dac_3v_8bit_0/b0a a_30098_n16820# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2715 dvss a_n53983_n17697# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2716 a_23170_n2566# vdd a_22563_n2963# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2717 dac_3v_column_0[7].res1_in vdd a_20863_n18713# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2718 dac_3v_column_odd_0[1].out_3 dac_3v_8bit_0/b3a dac_3v_column_odd_0[1].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2719 a_30098_n7227# a_31605_n7227# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2720 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2721 a_34426_n11252# vss a_34426_n11252# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2722 dac_3v_column_odd_0[2].out_5 dac_3v_8bit_0/b5a dac_3v_column_odd_0[2].out4 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2723 a_n40589_11447# bias_0.bi__pmirr_0.gate sbamuxm4_0/ibp[1] dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X2724 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2725 a_20156_n8962# vdd dac_3v_column_odd_0[2].dum_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2726 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2727 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2728 dvss level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b1a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2729 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2730 a_28398_n17214# dac_3v_8bit_0/b0a dac_3v_column_odd_0[6].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2731 a_20156_n17490# vdd a_20156_n17490# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2732 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2733 dvss level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b2a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2734 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2735 dac_3v_column_odd_0[7].dum_in0 vss a_34426_n19780# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2736 a_23877_n17214# dac_3v_8bit_0/b0a dac_3v_column_odd_0[6].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2737 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2738 a_n55599_n18241# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n55681_n18241# dvss sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2739 a_22174_2206# a_22174_2371# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X2740 a_24677_n20686# vdd a_24070_n21083# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2741 dac_3v_column_odd_0[6].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[6].res_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X2742 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2743 dac_3v_column_0[0].dum1_in dac_3v_column_0[0].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2744 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2745 dvss a_n53523_n22049# testbuffer_0.tb__mux_0.tbm__passgate_5.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2746 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C a_n55681_n22593# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2747 a_27636_2837# a_27998_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2748 a_20863_n5921# vss a_20863_n5921# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2749 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2750 dac_3v_column_0[5].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_0[5].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2751 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2752 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2753 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2754 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2755 a_20156_n13226# vss dac_3v_column_odd_0[4].dum_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2756 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2757 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2758 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2759 dac_3v_8bit_0/b0b level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2760 a_28398_n16147# a_29905_n16147# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2761 dac_3v_column_0[2].out1_0_1 dac_3v_8bit_0/b0b a_25577_n8292# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2762 dac_3v_column_0[0].out1_0_0 dac_3v_8bit_0/b0b a_22563_n4028# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2763 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2764 a_n32750_2575# a_n31275_1643# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X2765 dac_3v_column_odd_0[1].out1_0_1 dac_3v_8bit_0/b0a a_25577_n7227# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2766 a_27058_3107# b4 dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X2767 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2768 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2769 sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X2770 dac_3v_column_odd_0[6].res_out1 dac_3v_8bit_0/b0b dac_3v_column_0[7].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2771 a_22370_n16147# dac_3v_8bit_0/b0a dac_3v_column_0[6].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2772 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2773 dvdd testbuffer_0.tb__mux_0.tbm__passgate_1.en a_n48623_n15278# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X2774 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2775 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2776 dac_3v_column_odd_0[7].dum_in1 dac_3v_column_odd_0[7].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2777 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2778 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2779 dvss level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b6b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2780 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2781 a_20156_n5763# vdd dac_3v_column_0[1].dum1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2782 dac_3v_column_0[3].out1_0_1 dac_3v_8bit_0/b0a a_25577_n10424# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2783 a_28398_n7619# a_29905_n7619# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2784 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2785 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2786 a_20156_n4698# vss dac_3v_column_odd_0[0].dum_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2787 a_33719_n17490# vdd dac_3v_column_odd_0[6].res_out1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2788 dvdd testbuffer_0.tb__mux_0.tbm__passgate_4.en a_n47185_n21248# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X2789 dvss a_23802_3107# a_24742_3404# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X2790 dac_3v_column_0[7].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_0[7].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2791 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2792 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C a_n55681_n22593# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2793 dac_3v_column_0[7].out0_1_1 dac_3v_8bit_0/b2a dac_3v_column_0[7].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2794 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2795 dac_3v_column_0[5].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[5].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2796 a_n53523_n22049# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._17_.X dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2797 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2798 dac_3v_column_odd_0[1].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[1].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2799 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2800 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2801 dac_3v_8bit_0/b6b level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2802 sbamuxm4_0/vb[5] a_n32029_8404# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X2803 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2804 a_32520_2837# a_31942_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=1e+06u
X2805 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2806 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n53615_n20961# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2807 dvss dac_3v_8bit_0/b3a dac_3v_8bit_0/b3b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2808 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2809 a_25384_n15082# dac_3v_8bit_0/b0b dac_3v_column_odd_0[5].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2810 dvss a_32882_3404# a_32520_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2811 a_26891_n5487# a_28398_n5487# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2812 a_28398_n5487# dac_3v_8bit_0/b0a dac_3v_column_0[1].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2813 dvss dvss dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X2814 dvss a_23802_3107# a_23802_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2815 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2816 level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2817 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2818 a_31412_n7619# dac_3v_column_odd_0[1].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2819 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2820 dvss a_n54221_n17179# testbuffer_0.tb__mux_0.tbm__passgate_1.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2821 vdd dac_3v_8bit_0/b1a dac_3v_8bit_0/b1b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2822 a_30098_n10424# a_31605_n10424# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2823 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2824 vdd a_22174_2206# level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X2825 vdd level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2826 dac_3v_8bit_0/b0b level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2827 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2828 dac_3v_column_odd_0[3].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[3].res_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X2829 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2830 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2831 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2832 dac_3v_column_0[6].dum1_in dac_3v_column_0[6].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2833 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2834 dac_3v_8bit_0/b1b dac_3v_8bit_0/b1a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2835 dvss dac_3v_8bit_0/b0b dac_3v_8bit_0/b0a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2836 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2837 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2838 a_30705_n2566# vss a_30705_n2566# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2839 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output4.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n53825_n18785# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2840 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2841 dac_3v_column_odd_0[6].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[6].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2842 dac_3v_column_odd_0[5].out0_2 dac_3v_8bit_0/b3a dac_3v_column_odd_0[5].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2843 dac_3v_column_odd_0[7].in_5 vss dac_3v_column_odd_0[7].in_5 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=500000u
X2844 dac_3v_column_0[6].res1_in a_22563_n16820# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2845 dac_3v_8bit_0/b1b dac_3v_8bit_0/b1a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2846 a_22370_n7619# a_23877_n7619# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2847 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2848 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2849 a_23877_n18279# a_25384_n18279# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2850 a_22370_n2290# vdd a_22370_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2851 dac_3v_8bit_0/b3b dac_3v_8bit_0/b3a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2852 a_28591_n5095# a_30098_n5095# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2853 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2854 a_26891_n3355# dac_3v_8bit_0/b0a dac_3v_column_0[0].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2855 a_31412_n5487# dac_3v_8bit_0/b0a dac_3v_column_0[1].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2856 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2857 vdd level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b4a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2858 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2859 level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X2860 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2861 dvss bias_0.bi__amplifier_0.bias bias_0.bi__amplifier_0.bias dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X2862 dac_3v_column_0[3].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_0[3].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2863 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2864 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2865 dac_3v_column_odd_0[7].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[7].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2866 a_25577_n21083# a_27084_n21083# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2867 a_20863_n10185# vss a_20863_n10185# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2868 dac_3v_column_0[4].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_0[4].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2869 dvdd bias_0.bi__amplifier_0.mirr bias_0.bi__amplifier_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X2870 bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X2871 a_25384_n11883# dac_3v_8bit_0/b0b dac_3v_column_0[4].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2872 a_23170_n10818# dac_3v_8bit_0/b2b dac_3v_column_odd_0[3].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2873 dac_3v_column_odd_0[0].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_odd_0[0].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2874 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2875 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2876 dvdd a_n53615_n20961# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2877 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2878 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2879 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/muxout dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X2880 dac_3v_column_odd_0[0].res_in1 vdd a_20863_n4856# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2881 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2882 a_31605_n5095# dac_3v_column_odd_0[0].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2883 dac_3v_column_odd_0[5].res_in1 vdd a_20863_n15516# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2884 a_23170_n17214# dac_3v_8bit_0/b1a dac_3v_column_odd_0[6].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2885 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2886 dac_3v_column_0[7].out1_0_0 dac_3v_8bit_0/b0a a_22563_n18952# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2887 dac_3v_column_0[4].out1_0_2 dac_3v_8bit_0/b0a a_27084_n12556# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2888 dac_3v_column_0[0].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[0].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2889 dac_3v_column_0[4].out0_2 dac_3v_8bit_0/b3a dac_3v_column_0[4].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2890 dvss a_28686_3107# a_29626_3404# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X2891 dac_3v_column_odd_0[0].out_5 dac_3v_8bit_0/b6b dac_3v_column_odd_0[2].in_5 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2892 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2893 dac_3v_column_0[7].out_3 dac_3v_8bit_0/b3a dac_3v_column_0[7].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2894 a_26184_n2566# vss a_26184_n2566# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2895 dac_3v_column_odd_0[2].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_odd_0[2].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2896 dac_3v_column_odd_0[2].dum_out1 vss a_34426_n10185# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2897 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2898 a_n40589_12567# bias_0.bi__pmirr_0.gate sbamuxm4_0/ibp[3] dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X2899 a_23170_n20686# vdd a_23170_n20686# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2900 a_24070_n2963# a_25577_n2963# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2901 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2902 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n48623_n24233# inp[6] dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2903 a_22563_n5095# a_24070_n5095# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2904 a_26891_n20410# vss a_26891_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2905 vdd level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b5a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2906 dac_3v_column_odd_0[0].out_3 dac_3v_8bit_0/b3b dac_3v_column_odd_0[0].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2907 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2908 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2909 dac_3v_8bit_0/b4a level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2910 a_33719_n17490# vss dac_3v_column_odd_0[6].res_out1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X2911 dac_3v_column_odd_0[3].out4 dac_3v_8bit_0/b4b dac_3v_column_0[3].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2912 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2913 a_22563_n14688# a_24070_n14688# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2914 dac_3v_column_odd_0[2].dum_in1 dac_3v_column_odd_0[2].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2915 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2916 dac_3v_column_0[7].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_0[7].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2917 dac_3v_column_0[5].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[5].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2918 a_25384_n9751# dac_3v_8bit_0/b0b dac_3v_column_0[3].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2919 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2920 a_28398_n12950# a_29905_n12950# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2921 dac_3v_column_odd_0[0].out1_0_2 dac_3v_8bit_0/b0b a_27084_n5095# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2922 dvdd a_n55646_9265# bias_basis_current_0.bb__pmirr_0.vbn dvss sky130_fd_pr__nfet_01v8_lvt ad=2.22214e+14p pd=2.56439e+09u as=0p ps=0u w=1e+06u l=300000u
X2923 a_29905_n20844# vss a_29905_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2924 dac_3v_column_odd_0[2].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_odd_0[2].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2925 a_26891_n14015# a_28398_n14015# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2926 bias_0.bi__amplifier_0.bias bias_0.bi__amplifier_0.bias dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X2927 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2928 dac_3v_column_0[6].out1_0_1 dac_3v_8bit_0/b0b a_24070_n16820# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2929 dac_3v_column_odd_0[5].res_in0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[5].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2930 dac_3v_column_0[2].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[2].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2931 vdd level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2932 level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2933 dac_3v_column_0[3].out1_0_2 dac_3v_8bit_0/b0b a_28591_n10424# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2934 dac_3v_column_odd_0[1].out1_0_3 dac_3v_8bit_0/b0b a_31605_n7227# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X2935 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2936 dac_3v_column_0[4].res1_in vdd a_20863_n12317# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2937 dac_3v_8bit_0/b5a level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2938 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output6.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2939 a_24070_n6160# a_25577_n6160# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2940 dac_3v_column_odd_0[5].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_odd_0[5].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2941 a_26891_n16147# dac_3v_8bit_0/b0b dac_3v_column_0[6].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2942 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2943 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2944 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2945 a_25577_n9359# a_27084_n9359# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2946 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X2947 dac_3v_column_0[1].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_0[1].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2948 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2949 a_22370_n16147# dac_3v_8bit_0/b0b dac_3v_column_0[6].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2950 dac_3v_column_odd_0[2].out4 dac_3v_8bit_0/b4a dac_3v_column_0[2].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2951 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2952 dac_3v_8bit_0/b5b dac_3v_8bit_0/b5a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2953 a_20863_n20410# a_22370_n20410# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2954 dac_3v_column_odd_0[2].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[2].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2955 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X2956 dac_3v_column_odd_0[4].res_out1 dac_3v_column_odd_0[4].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2957 a_29905_n9751# dac_3v_8bit_0/b0a dac_3v_column_0[3].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X2958 dac_3v_column_0[1].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[1].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X2959 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2960 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbn dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2961 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2962 dac_3v_column_odd_0[5].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_odd_0[5].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2963 a_23170_n15082# dac_3v_8bit_0/b2a dac_3v_column_odd_0[5].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2964 a_33719_n7895# vdd dac_3v_column_odd_0[2].res_in0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X2965 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2966 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2967 a_24070_n12556# a_25577_n12556# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2968 a_23170_n8686# dac_3v_8bit_0/b2a dac_3v_column_odd_0[2].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X2969 a_n46909_n18263# a_n47185_n18263# dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X2970 dac_3v_column_odd_0[5].out1_0_2 dac_3v_8bit_0/b0b a_27084_n15755# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2971 dac_3v_column_0[2].dum1_in dac_3v_column_0[2].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2972 dac_3v_column_0[2].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[2].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2973 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2974 level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=2.1e+11p pd=2.06e+06u as=0p ps=0u w=750000u l=500000u
X2975 dac_3v_column_0[2].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[2].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X2976 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X2977 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X2978 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2979 a_n26631_n925# a_n26245_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X2980 a_28686_2371# a_29264_2837# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.142e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=1e+06u
X2981 a_14987_n11444# a_14987_n11444# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2982 dac_3v_column_odd_0[7].out1_0_3 dac_3v_8bit_0/b0a a_31605_n20019# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2983 dvdd a_n55547_n19873# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2984 a_n54345_n20265# a_n54072_n20437# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2985 a_n54691_n21255# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n54945_n21255# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2986 a_26891_n2290# a_28398_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2987 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X2988 a_30098_n4028# a_31605_n4028# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X2989 dac_3v_column_0[2].out1_0_1 dac_3v_8bit_0/b0b a_24070_n8292# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2990 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2991 dac_3v_column_0[1].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_0[1].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X2992 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2993 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2994 dac_3v_column_odd_0[3].res_out1 dac_3v_8bit_0/b0b dac_3v_column_0[4].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X2995 dvss a_31254_3404# a_30892_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2996 dac_3v_column_0[2].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[2].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2997 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2998 a_28398_n14015# dac_3v_8bit_0/b0a dac_3v_column_0[5].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X2999 a_20156_n14291# vdd a_20156_n14291# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3000 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3001 a_29905_n15082# a_31412_n15082# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3002 dac_3v_column_odd_0[4].dum_in1 dac_3v_column_odd_0[4].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3003 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3004 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3005 dac_3v_column_odd_0[5].dum_out1 vss a_34426_n16581# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3006 a_23877_n14015# dac_3v_8bit_0/b0a dac_3v_column_0[5].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3007 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3008 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3009 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3010 a_23802_2371# a_23802_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3011 a_31605_n15755# dac_3v_column_odd_0[5].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3012 dac_3v_column_odd_0[4].res_in1 a_22563_n13623# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3013 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3014 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3015 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3016 dac_3v_column_0[1].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_0[1].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3017 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3018 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X3019 dac_3v_column_0[5].out1_0_1 dac_3v_8bit_0/b0a a_25577_n14688# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3020 a_20156_n10027# vss dac_3v_column_0[3].dum1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3021 a_34426_n18713# vdd a_34426_n18713# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3022 vdd level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b0b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3023 dac_3v_column_0[4].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_0[4].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3024 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3025 a_n54482_n20601# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n54563_n20601# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.071e+11p ps=1.35e+06u w=420000u l=150000u
X3026 level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3027 a_20863_n15516# vdd a_20863_n15516# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3028 dac_3v_column_0[4].out0_1_1 dac_3v_8bit_0/b2a dac_3v_column_0[4].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3029 dac_3v_8bit_0/b0a dac_3v_8bit_0/b0b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3030 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3031 dac_3v_column_0[2].out1_0_2 dac_3v_8bit_0/b0a a_27084_n8292# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3032 a_29905_n6554# dac_3v_8bit_0/b0b dac_3v_column_odd_0[1].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3033 dac_3v_column_0[0].out1_0_1 dac_3v_8bit_0/b0a a_24070_n4028# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3034 vdd level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
D7 dvss b7 sky130_fd_pr__diode_pw2nd_05v5
X3035 dac_3v_column_odd_0[7].dum_out1 vdd a_34426_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3036 a_23170_n12950# dac_3v_8bit_0/b1b dac_3v_column_odd_0[4].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3037 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3038 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3039 a_26891_n12950# dac_3v_8bit_0/b0a dac_3v_column_odd_0[4].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X3040 dvdd bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbp dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3041 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3042 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n53615_n20961# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3043 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3044 bandgap_0.bg__pnp_group_0.eg dvss a_n31275_2703# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X3045 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3046 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3047 bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3048 a_n54937_n18785# a_n55047_n18669# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output6.A dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3049 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X3050 dac_3v_column_0[7].out1_0_1 dac_3v_8bit_0/b0b a_25577_n18952# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3051 a_31412_n17214# dac_3v_8bit_0/b0b dac_3v_column_odd_0[6].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3052 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3053 dvdd w_n19679_n3822# a_n21740_n3691# dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X3054 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X3055 dvss dac_3v_8bit_0/b7b dac_3v_8bit_0/b7a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3056 dvss level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b3a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3057 a_32212_n20686# vdd a_31605_n21083# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3058 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3059 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3060 dvss a_n54301_n18241# testbuffer_0.tb__mux_0.tbm__passgate_3.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3061 a_31942_3107# b1 dvss dvss sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X3062 a_28591_n17887# a_30098_n17887# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3063 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3064 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._19_.A a_n54487_n21933# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3065 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3066 dac_3v_column_odd_0[0].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[0].res_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3067 dac_3v_column_odd_0[7].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_odd_0[7].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3068 a_26184_n20686# vss a_26184_n20686# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3069 a_29905_n10818# dac_3v_8bit_0/b0a dac_3v_column_odd_0[3].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3070 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3071 dac_3v_column_odd_0[0].res_in0 dac_3v_column_odd_0[0].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3072 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3073 dac_3v_column_odd_0[1].dum_in0 vdd a_34426_n6988# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X3074 dvss dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inn sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=1
X3075 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3076 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3077 dac_3v_column_0[0].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[0].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3078 dac_3v_column_odd_0[6].out0_2 dac_3v_8bit_0/b3b dac_3v_column_odd_0[6].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X3079 dac_3v_column_odd_0[5].out4 dac_3v_8bit_0/b4b dac_3v_column_odd_0[5].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3080 dac_3v_column_odd_0[4].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[4].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3081 dvss level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b7b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3082 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3083 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3084 dac_3v_column_odd_0[3].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_odd_0[3].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3085 a_n32750_n4845# a_n31275_n4717# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X3086 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3087 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3088 dvss a_n55353_n19355# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3089 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3090 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3091 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/muxout dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X3092 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3093 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3094 a_28398_n19346# dac_3v_8bit_0/b0b dac_3v_column_odd_0[7].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3095 a_22563_n11491# a_24070_n11491# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3096 a_25384_n6554# dac_3v_8bit_0/b0a dac_3v_column_odd_0[1].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3097 a_n42353_11671# bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3098 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3099 dac_3v_column_odd_0[5].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_odd_0[5].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3100 dvss a_33570_2206# level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X3101 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3102 dac_3v_column_0[5].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_0[5].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X3103 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3104 a_32919_n2290# vdd a_32919_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X3105 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3106 dac_3v_column_odd_0[5].out1_0_3 dac_3v_8bit_0/b0b a_30098_n15755# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3107 a_20863_n14449# vss a_20863_n14449# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3108 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3109 dac_3v_column_odd_0[5].out1_0_1 dac_3v_8bit_0/b0a a_24070_n15755# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3110 dvdd bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbp dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3111 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3112 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X3113 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
D8 dvss b0 sky130_fd_pr__diode_pw2nd_05v5
X3114 dac_3v_column_odd_0[0].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[0].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3115 dac_3v_column_odd_0[6].out_5 dac_3v_8bit_0/b5b dac_3v_column_odd_0[6].out4 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3116 a_26891_n10818# a_28398_n10818# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3117 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3118 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3119 dac_3v_8bit_0/b4a level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3120 a_33719_n2566# vdd a_33719_n2566# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3121 a_16155_n11444# a_16155_n11444# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X3122 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3123 a_11923_n7894# a_17355_n8212# vss sky130_fd_pr__res_xhigh_po w=350000u l=2.5e+07u
X3124 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3125 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3126 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3127 dac_3v_8bit_0/b5b dac_3v_8bit_0/b5a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3128 a_33719_n8962# vss dac_3v_column_odd_0[2].res_out1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3129 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3130 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3131 a_23877_n2290# vdd a_23877_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3132 a_28398_n2724# vdd a_28398_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3133 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3134 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3135 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3136 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3137 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3138 a_31412_n20844# vdd a_31412_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3139 dac_3v_column_odd_0[6].dum_in1 dac_3v_column_odd_0[6].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3140 a_24070_n20019# a_25577_n20019# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3141 dac_3v_column_0[6].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[6].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3142 dac_3v_column_odd_0[3].res_in0 dac_3v_column_odd_0[3].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3143 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3144 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3145 bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas bias_0.bi__pmirr_0.gate_cas dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3146 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3147 dvss dac_3v_8bit_0/b7b dac_3v_8bit_0/b7a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3148 a_24677_n2566# vdd a_24677_n2566# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3149 sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X3150 dvdd bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3151 dac_3v_column_odd_0[2].res_in0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[2].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3152 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3153 vdd a_16155_n11444# follower_amp_0.pdrv2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3154 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3155 dac_3v_column_0[3].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_0[3].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3156 vdd level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3157 dac_3v_column_odd_0[0].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[0].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3158 a_n54563_n20601# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3159 dac_3v_column_0[7].out0_1_1 dac_3v_8bit_0/b2b dac_3v_column_0[7].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3160 a_n32750_455# a_n31275_583# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X3161 dac_3v_8bit_0/b1a level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3162 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3163 bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X3164 a_23877_n17214# a_25384_n17214# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3165 dac_3v_column_odd_0[5].out4 dac_3v_8bit_0/b4b dac_3v_column_0[5].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3166 dac_3v_column_0[4].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_0[4].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3167 dac_3v_column_odd_0[3].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[3].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3168 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3169 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3170 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X3171 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3172 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3173 a_30314_2371# a_30892_2837# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.142e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=1e+06u
X3174 a_22370_n9751# dac_3v_8bit_0/b0a dac_3v_column_0[3].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3175 dac_3v_column_0[5].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[5].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3176 dac_3v_column_0[3].res1_in a_22370_n9751# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3177 a_31412_n2724# vdd a_31412_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3178 a_31412_n18279# dac_3v_column_odd_0[6].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3179 dac_3v_column_odd_0[4].dum_in0 vdd a_34426_n13384# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3180 a_23877_n19346# dac_3v_8bit_0/b0b dac_3v_column_odd_0[7].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3181 a_23877_n8686# dac_3v_8bit_0/b0a dac_3v_column_odd_0[2].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3182 dac_3v_column_odd_0[1].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[1].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3183 dac_3v_8bit_0/b7a dac_3v_8bit_0/b7b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3184 a_23170_n4422# dac_3v_8bit_0/b1b dac_3v_column_odd_0[0].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3185 a_29905_n8686# a_31412_n8686# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3186 a_27691_n2566# vss a_27691_n2566# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3187 dac_3v_column_0[7].out1_0_3 dac_3v_8bit_0/b0b a_31605_n18952# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3188 dac_3v_column_0[5].out1_0_2 dac_3v_8bit_0/b0b a_28591_n14688# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3189 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3190 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3191 a_33719_n5763# vss dac_3v_column_odd_0[1].res_in0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3192 a_n41084_7938# bias_0.bi__nmirr_0.gate_n dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X3193 dac_3v_8bit_0/b7a dac_3v_8bit_0/b7b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3194 dac_3v_column_odd_0[3].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[3].res_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3195 a_25577_n2963# a_27084_n2963# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3196 dac_3v_column_odd_0[2].out1_0_2 dac_3v_8bit_0/b0b a_28591_n9359# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3197 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3198 dac_3v_column_odd_0[3].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[3].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3199 a_32212_n20686# vss a_32212_n20686# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3200 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._19_.X a_n53197_n22593# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3201 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3202 a_30892_2837# a_31254_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3203 dac_3v_column_0[1].dum1_in dac_3v_column_0[1].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3204 dac_3v_column_odd_0[7].in_5 vdd dac_3v_column_odd_0[7].in_5 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X3205 a_23170_n12950# dac_3v_8bit_0/b1b dac_3v_column_odd_0[4].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3206 dvss testbuffer_0.tb__mux_0.tbm__passgate_0.en a_n47185_n15278# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X3207 sbamuxm4_0/ibp[0] sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3208 dvdd a_30314_3107# a_31254_3404# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X3209 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3210 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3211 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3212 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3213 dac_3v_column_odd_0[0].out4 dac_3v_8bit_0/b4b dac_3v_column_0[0].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3214 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3215 sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X3216 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n53553_n18785# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3217 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3218 a_34426_n6988# vdd a_34426_n6988# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3219 dac_3v_column_0[3].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[3].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3220 a_n47950_6120# bias_0.bi__amplifier_0.bias bias_0.bi__amplifier_0.diff dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X3221 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out bias_0.bi__amplifier_0.inn dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3222 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3223 w_n19679_n3822# dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3224 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X3225 dvss level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3226 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3227 dac_3v_column_0[4].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_0[4].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3228 a_n23543_n925# a_n24315_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X3229 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3230 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3231 dvss level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3232 a_25577_n6160# a_27084_n6160# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3233 dac_3v_column_0[2].out_3 dac_3v_8bit_0/b3a dac_3v_column_0[2].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3234 dac_3v_column_0[0].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[0].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X3235 dac_3v_column_odd_0[1].res_in1 a_22563_n7227# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3236 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3237 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3238 a_30098_n8292# a_31605_n8292# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3239 dac_3v_column_odd_0[1].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_odd_0[1].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3240 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3241 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3242 dac_3v_column_odd_0[5].out1_0_3 dac_3v_8bit_0/b0a a_30098_n15755# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3243 a_33719_n11094# vdd dac_3v_column_odd_0[3].res_out1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3244 dvss bias_0.bi__nmirr_0.gate_n dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3245 dac_3v_column_0[1].out0_1_1 dac_3v_8bit_0/b2a dac_3v_column_0[1].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X3246 dac_3v_column_0[1].out1_0_2 dac_3v_8bit_0/b0b a_28591_n6160# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3247 a_20156_n6830# vss a_20156_n6830# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X3248 a_33719_n19622# vdd a_33719_n19622# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3249 dac_3v_column_0[4].out1_0_2 dac_3v_8bit_0/b0b a_27084_n12556# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3250 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3251 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inp bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3252 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3253 vdd dac_3v_8bit_0/b4a dac_3v_8bit_0/b4b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3254 dac_3v_8bit_0/b0a dac_3v_8bit_0/b0b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3255 dac_3v_column_0[6].out1_0_3 dac_3v_8bit_0/b0a a_31605_n16820# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3256 a_20156_n14291# vss dac_3v_column_0[5].dum1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3257 a_20863_n4856# vss a_20863_n4856# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3258 dac_3v_column_odd_0[4].out_3 dac_3v_8bit_0/b3b dac_3v_column_odd_0[4].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X3259 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3260 dac_3v_column_odd_0[4].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[4].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3261 a_31412_n10818# dac_3v_8bit_0/b0a dac_3v_column_odd_0[3].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3262 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3263 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3264 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3265 sbamuxm4_0/ibn[0] bias_0.bi__pmirr_0.gate_cas a_n41084_8994# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3266 dac_3v_column_0[2].out1_0_1 dac_3v_8bit_0/b0a a_25577_n8292# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3267 a_n41084_7586# bias_0.bi__nmirr_0.gate_n dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3268 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3269 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3270 a_23170_n2566# vss a_22563_n2963# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3271 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3272 a_29905_n11883# a_31412_n11883# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3273 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3274 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3275 dac_3v_column_odd_0[3].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[3].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3276 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3277 dac_3v_8bit_0/b3b dac_3v_8bit_0/b3a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3278 dac_3v_column_0[3].res1_in a_22563_n10424# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3279 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inp bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
D9 dvss b2 sky130_fd_pr__diode_pw2nd_05v5
X3280 a_31605_n12556# dac_3v_column_odd_0[4].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3281 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3282 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3283 a_29905_n19346# dac_3v_8bit_0/b0b dac_3v_column_odd_0[7].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3284 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3285 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3286 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3287 dac_3v_column_0[7].out1_0_2 dac_3v_8bit_0/b0a a_28591_n18952# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3288 a_20863_n12317# vdd a_20863_n12317# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3289 a_n54657_n18785# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3290 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3291 a_29905_n3355# dac_3v_8bit_0/b0b dac_3v_column_0[0].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3292 a_20156_n4698# vdd dac_3v_column_odd_0[0].dum_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3293 testbuffer_0.tb__mux_0.tbm__passgate_5.en a_n53523_n22049# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3294 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3295 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3296 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3297 a_28686_2371# a_28686_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3298 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3299 a_29198_n20686# vdd a_29198_n20686# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3300 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3301 a_27084_n18952# a_28591_n18952# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3302 a_34426_n13384# vss a_34426_n13384# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3303 dac_3v_8bit_0/b5a level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3304 dac_3v_column_odd_0[4].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[4].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3305 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3306 a_23170_n15082# dac_3v_8bit_0/b2b dac_3v_column_odd_0[5].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3307 a_31412_n14015# dac_3v_8bit_0/b0b dac_3v_column_0[5].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3308 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3309 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3310 a_28591_n14688# a_30098_n14688# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3311 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3312 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3313 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3314 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3315 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3316 dac_3v_column_0[6].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_0[6].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3317 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3318 dac_3v_column_odd_0[7].res_in0 dac_3v_column_odd_0[7].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3319 dac_3v_column_0[0].dum0_in vdd a_34426_n3789# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3320 dac_3v_column_odd_0[7].out1_0_1 dac_3v_8bit_0/b0a a_25577_n20019# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3321 a_29905_n18279# dac_3v_8bit_0/b0a dac_3v_column_0[7].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3322 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3323 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3324 dac_3v_column_0[5].out0_2 dac_3v_8bit_0/b3b dac_3v_column_0[5].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X3325 dac_3v_column_odd_0[4].out4 dac_3v_8bit_0/b4a dac_3v_column_0[4].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3326 dac_3v_column_0[3].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_0[3].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3327 dvss a_33570_3107# a_33570_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3328 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3329 dvss bias_0.bi__nmirr_0.gate_n bias_0.bi__nmirr_0.gate_n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3330 a_22752_2837# a_22174_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=1e+06u
X3331 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3332 dvss a_n53523_n22049# testbuffer_0.tb__mux_0.tbm__passgate_5.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3333 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3334 a_33719_n11094# vss dac_3v_column_odd_0[3].res_out1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X3335 dvss dac_3v_8bit_0/b2a dac_3v_8bit_0/b2b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3336 a_25384_n3355# dac_3v_8bit_0/b0a dac_3v_column_0[0].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3337 a_28398_n16147# dac_3v_8bit_0/b0b dac_3v_column_0[6].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3338 vdd dac_3v_8bit_0/b7b dac_3v_8bit_0/b7a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3339 a_20024_n2963# a_20863_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3340 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3341 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3342 a_n42353_12119# bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3343 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X3344 a_26891_n6554# dac_3v_8bit_0/b0b dac_3v_column_odd_0[1].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3345 a_26891_n2290# vss a_26891_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3346 a_33719_n19622# vss a_33719_n19622# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3347 a_25577_n15755# a_27084_n15755# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3348 a_n48347_n21248# a_n48623_n21248# dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X3349 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3350 dac_3v_column_0[4].out1_0_3 dac_3v_8bit_0/b0b a_30098_n12556# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3351 a_20156_n18555# vdd dac_3v_column_0[7].dum1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3352 dac_3v_column_0[7].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_0[7].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3353 dac_3v_column_0[4].out1_0_1 dac_3v_8bit_0/b0a a_24070_n12556# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3354 a_28398_n9751# a_29905_n9751# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3355 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3356 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3357 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3358 dac_3v_column_0[7].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[7].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3359 dac_3v_column_0[4].out0_1_1 dac_3v_8bit_0/b2b dac_3v_column_0[4].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3360 a_20156_n6830# vss dac_3v_column_odd_0[1].dum_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3361 vdd dac_3v_8bit_0/b5a dac_3v_8bit_0/b5b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3362 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3363 dac_3v_column_odd_0[1].out0_2 dac_3v_8bit_0/b3a dac_3v_column_odd_0[1].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3364 level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X3365 w_n19679_n3822# dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3366 dvss level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b2a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3367 a_20156_n20686# vdd a_20156_n20686# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3368 a_28398_n20410# vdd a_28398_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3369 level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3370 vdd level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b6b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3371 sbamuxm4_0/ibn[1] bias_0.bi__pmirr_0.gate_cas a_n41084_9346# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3372 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3373 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3374 a_23877_n20410# vss a_23877_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3375 dvss a_22174_2206# level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X3376 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3377 dac_3v_8bit_0/b5a level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3378 dac_3v_column_0[5].dum1_in dac_3v_column_0[5].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3379 a_25384_n17214# dac_3v_8bit_0/b0b dac_3v_column_odd_0[6].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3380 dac_3v_column_odd_0[6].out1_0_0 dac_3v_8bit_0/b0a a_22563_n17887# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3381 a_26184_n20686# vdd a_25577_n21083# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3382 a_28398_n7619# dac_3v_8bit_0/b0a dac_3v_column_0[2].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3383 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3384 dac_3v_column_odd_0[2].res_out1 dac_3v_8bit_0/b0b dac_3v_column_0[3].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3385 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3386 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3387 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n47185_n15278# inp[0] dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3388 a_26184_n2566# vdd a_26184_n2566# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3389 dac_3v_column_odd_0[0].res_out1 dac_3v_8bit_0/b0a dac_3v_column_0[1].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=500000u
X3390 dac_3v_column_odd_0[6].out_3 dac_3v_8bit_0/b3a dac_3v_column_odd_0[6].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3391 a_31412_n9751# dac_3v_column_odd_0[2].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3392 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3393 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3394 a_28686_3107# b3 dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X3395 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3396 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3397 dac_3v_column_odd_0[7].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_odd_0[7].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3398 dac_3v_column_odd_0[4].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[4].res_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3399 dac_3v_column_odd_0[2].dum_in0 vss a_34426_n9120# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3400 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3401 a_20863_n19780# vss a_20863_n19780# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3402 a_23877_n14015# a_25384_n14015# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3403 a_33719_n10027# vdd a_33719_n10027# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X3404 dvss bias_0.bi__pmirr_0.gate_cas dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3405 a_25430_3107# b5 dvss dvss sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X3406 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3407 a_34148_2837# a_33570_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=1e+06u
X3408 dac_3v_8bit_0/b3a level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3409 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3410 bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X3411 dac_3v_8bit_0/b0a dac_3v_8bit_0/b0b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3412 dac_3v_column_odd_0[6].out0_2 dac_3v_8bit_0/b3a dac_3v_column_odd_0[6].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X3413 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inn bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3414 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3415 a_23877_n9751# dac_3v_8bit_0/b0b dac_3v_column_0[3].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3416 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3417 w_n19679_n3822# dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3418 a_23877_n16147# dac_3v_8bit_0/b0b dac_3v_column_0[6].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3419 a_22370_n9751# a_23877_n9751# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3420 a_31942_2371# a_32520_2837# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.142e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=1e+06u
X3421 a_23877_n5487# dac_3v_8bit_0/b0a dac_3v_column_0[1].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3422 dvss bias_0.bi__nmirr_0.gate_n bias_0.bi__nmirr_0.gate_n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3423 dvss a_n54441_n21531# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output8.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3424 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._19_.A a_n53289_n21505# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3425 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3426 dac_3v_column_odd_0[4].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[4].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3427 a_25384_n8686# dac_3v_8bit_0/b0b dac_3v_column_odd_0[2].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X3428 a_28591_n7227# a_30098_n7227# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3429 a_29905_n5487# a_31412_n5487# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3430 a_31412_n7619# dac_3v_8bit_0/b0a dac_3v_column_0[2].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3431 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3432 dac_3v_column_0[3].out0_1_1 dac_3v_8bit_0/b2b dac_3v_column_0[3].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3433 dac_3v_column_0[2].out1_0_3 dac_3v_8bit_0/b0b a_31605_n8292# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3434 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3435 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3436 dac_3v_8bit_0/b5a level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3437 a_31605_n20019# vlow vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3438 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X3439 dvss a_25430_3107# a_25430_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3440 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3441 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3442 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3443 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3444 dac_3v_column_odd_0[5].out1_0_1 dac_3v_8bit_0/b0b a_24070_n15755# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3445 dac_3v_column_odd_0[2].out1_0_3 dac_3v_8bit_0/b0b a_30098_n9359# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3446 a_n21999_n925# a_n20841_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X3447 dvss a_n53615_n20961# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3448 dac_3v_column_odd_0[6].out_5 dac_3v_8bit_0/b5a dac_3v_column_odd_0[6].out4 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3449 vdd a_16155_n11444# a_16155_n11444# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3450 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3451 dac_3v_column_0[7].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[7].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3452 dac_3v_column_odd_0[5].res_in1 a_22370_n15082# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3453 a_31412_n17214# dac_3v_column_odd_0[6].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3454 bias_0.bi__amplifier_0.mirr bias_0.bi__pmirr_0.fb bias_0.bi__amplifier_0.diff dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X3455 a_20863_n9120# vdd a_20863_n9120# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3456 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3457 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3458 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3459 dac_3v_column_odd_0[0].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_odd_0[0].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3460 a_26891_n19346# a_28398_n19346# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3461 dac_3v_column_odd_0[7].out4 dac_3v_8bit_0/b4a dac_3v_column_odd_0[7].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3462 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3463 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3464 dvdd a_31942_3107# a_32882_3404# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X3465 level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3466 vdd dac_3v_8bit_0/b3a dac_3v_8bit_0/b3b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3467 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3468 a_34426_n3789# vss a_34426_n3789# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3469 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3470 dac_3v_column_odd_0[6].res_in1 vdd a_20863_n17648# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3471 a_31605_n7227# dac_3v_column_odd_0[1].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3472 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X3473 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3474 vdd level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3475 a_29905_n8686# dac_3v_8bit_0/b0a dac_3v_column_odd_0[2].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3476 dac_3v_column_odd_0[2].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[2].res_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3477 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output4.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3478 a_n46909_n21248# a_n47185_n21248# dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X3479 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3480 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3481 a_25384_n20844# vdd a_25384_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3482 dac_3v_column_0[3].out0_2 dac_3v_8bit_0/b3b dac_3v_column_0[3].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3483 bias_0.bi__amplifier_0.diff bias_0.bi__pmirr_0.fb bias_0.bi__amplifier_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X3484 a_20863_n20844# vss a_20863_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3485 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3486 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3487 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3488 dac_3v_column_odd_0[7].res_in0 dac_3v_column_odd_0[7].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3489 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3490 dac_3v_column_0[0].res1_in a_22563_n4028# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3491 dac_3v_column_odd_0[7].out1_0_2 dac_3v_8bit_0/b0b a_28591_n20019# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3492 a_28591_n11491# a_30098_n11491# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3493 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3494 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3495 dac_3v_8bit_0/b7b level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3496 dac_3v_column_0[4].out1_0_3 dac_3v_8bit_0/b0a a_30098_n12556# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3497 a_22563_n7227# a_24070_n7227# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3498 dvdd bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3499 dac_3v_column_0[0].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_0[0].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3500 dac_3v_column_odd_0[1].out_3 dac_3v_8bit_0/b3b dac_3v_column_odd_0[1].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3501 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output5.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3502 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3503 dac_3v_column_odd_0[0].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_odd_0[0].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3504 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3505 dvss level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3506 vdd level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b5a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3507 a_20156_n3631# vss a_20156_n3631# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3508 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3509 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3510 a_22563_n16820# a_24070_n16820# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3511 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X a_n53983_n17697# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3512 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3513 a_33719_n16423# vdd a_33719_n16423# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3514 a_29905_n15082# dac_3v_8bit_0/b0a dac_3v_column_odd_0[5].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3515 a_n47950_6120# bias_0.bi__amplifier_0.bias dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X3516 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3517 sbamuxm4_0/ibp[0] sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3518 dac_3v_column_0[1].out1_0_3 dac_3v_8bit_0/b0b a_30098_n6160# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3519 a_25384_n18279# a_26891_n18279# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3520 dac_3v_8bit_0/out_unbuf dac_3v_8bit_0/b7a dac_3v_column_odd_0[2].in_5 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3521 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3522 a_28398_n12950# dac_3v_8bit_0/b0a dac_3v_column_odd_0[4].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3523 a_20156_n13226# vdd a_20156_n13226# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3524 dac_3v_column_odd_0[1].out1_0_2 dac_3v_8bit_0/b0b a_27084_n7227# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3525 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3526 a_n46909_n24233# a_n47185_n24233# dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X3527 dac_3v_8bit_0/b1a level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3528 dvdd a_n55233_n20443# testbuffer_0.tb__mux_0.tbm__passgate_4.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3529 a_23877_n12950# dac_3v_8bit_0/b0a dac_3v_column_odd_0[4].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3530 sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X3531 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3532 dac_3v_8bit_0/b2b dac_3v_8bit_0/b2a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3533 dvss a_n54713_n20729# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._07_.X dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3534 a_20863_n5921# vdd a_20863_n5921# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3535 bias_0.bi__amplifier_0.diff bias_0.bi__pmirr_0.fb bias_0.bi__amplifier_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X3536 a_26891_n16147# a_28398_n16147# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3537 dac_3v_column_odd_0[6].res_in0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[6].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3538 dac_3v_column_0[3].out_3 dac_3v_8bit_0/b3b dac_3v_column_0[3].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X3539 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3540 dvss level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b0b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3541 dac_3v_column_odd_0[0].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[0].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3542 dac_3v_column_0[7].out1_0_0 dac_3v_8bit_0/b0b a_22563_n18952# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3543 a_n42000_8994# bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[0] dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X3544 dac_3v_column_0[3].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_0[3].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3545 a_34426_n17648# vdd a_34426_n17648# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3546 bias_0.bi__pmirr_0.fb a_n32029_12624# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X3547 dac_3v_column_0[1].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_0[1].res1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3548 a_32919_n20844# vss a_32919_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3549 a_23170_n10818# dac_3v_8bit_0/b1a dac_3v_column_odd_0[3].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=500000u
X3550 a_33570_2371# a_33570_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3551 dac_3v_8bit_0/b4b dac_3v_8bit_0/b4a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3552 dac_3v_column_0[0].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[0].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3553 a_31412_n18279# dac_3v_8bit_0/b0a dac_3v_column_0[7].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3554 bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inp a_n27403_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X3555 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3556 a_23170_n20686# vss a_23170_n20686# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3557 a_24677_n2566# vss a_24070_n2963# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3558 dac_3v_column_odd_0[5].res_out1 dac_3v_column_odd_0[5].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3559 a_n32750_n1665# a_n31275_n1537# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X3560 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3561 bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X3562 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3563 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3564 dac_3v_column_0[2].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[2].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3565 dac_3v_column_odd_0[6].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_odd_0[6].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3566 a_23170_n17214# dac_3v_8bit_0/b2a dac_3v_column_odd_0[6].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3567 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3568 a_29905_n16147# dac_3v_8bit_0/b0b dac_3v_column_0[6].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3569 vdd level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b4a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3570 dac_3v_column_odd_0[6].out1_0_1 dac_3v_8bit_0/b0b a_25577_n17887# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3571 a_29198_n20686# vss a_28591_n21083# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3572 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3573 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n48347_n15278# inp[1] dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3574 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3575 dvss a_28686_3107# a_28686_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3576 a_29905_n11883# dac_3v_8bit_0/b0a dac_3v_column_0[4].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3577 a_23877_n4422# a_25384_n4422# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3578 a_20156_n19622# vss dac_3v_column_odd_0[7].dum_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3579 dac_3v_column_odd_0[3].dum_in1 dac_3v_column_odd_0[3].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3580 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3581 bias_0.bi__amplifier_0.diff bias_0.bi__amplifier_0.bias a_n47950_6120# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X3582 level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3583 a_28398_n4422# dac_3v_8bit_0/b0a dac_3v_column_odd_0[0].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3584 a_n32750_n3785# a_n31275_n3657# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X3585 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3586 dac_3v_column_0[5].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_0[5].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3587 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3588 a_34426_n10185# vss a_34426_n10185# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3589 a_25430_3107# b5 dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X3590 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3591 a_32212_n2566# vss a_32212_n2566# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3592 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3593 a_23877_n10818# a_25384_n10818# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3594 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3595 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3596 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3597 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3598 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3599 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X3600 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3601 dac_3v_8bit_0/b4b dac_3v_8bit_0/b4a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3602 dac_3v_column_0[6].out1_0_1 dac_3v_8bit_0/b0a a_25577_n16820# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3603 bandgap_0.bg__se_folded_cascode_p_0.bgfc__diffpair_p_0.inp a_n31275_2703# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X3604 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3605 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3606 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._17_.X a_n55405_n20961# dvss dvss sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3607 dvdd a_n53615_n20961# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3608 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3609 a_29905_n2290# a_31412_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3610 a_31412_n4422# dac_3v_8bit_0/b0a dac_3v_column_odd_0[0].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3611 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3612 vdd level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b3a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3613 a_25384_n10818# dac_3v_8bit_0/b0a dac_3v_column_odd_0[3].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3614 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n46909_n18263# inp[3] dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3615 dac_3v_column_odd_0[3].res_in1 vss a_20863_n11252# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3616 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n54072_n20437# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.0785e+11p ps=1.36e+06u w=420000u l=150000u
X3617 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3618 a_22370_n20410# a_23877_n20410# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3619 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3620 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3621 a_25430_2206# a_25430_2371# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X3622 level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3623 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3624 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3625 a_n42353_11895# bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3626 dac_3v_column_odd_0[5].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[5].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3627 dvss level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3628 a_26891_n3355# dac_3v_8bit_0/b0b dac_3v_column_0[0].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3629 a_33719_n16423# vss a_33719_n16423# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3630 a_25577_n12556# a_27084_n12556# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3631 a_20156_n20686# vss a_20024_n21083# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3632 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3633 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3634 dvss a_22174_3107# a_22174_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3635 dvdd bias_0.bi__pmirr_0.gate a_n40589_11671# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3636 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3637 dac_3v_column_0[0].out0_2 dac_3v_8bit_0/b3a dac_3v_column_0[0].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3638 dac_3v_column_odd_0[5].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[5].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3639 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3640 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3641 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3642 dac_3v_column_odd_0[1].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[1].res_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=500000u
X3643 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3644 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3645 a_n42000_9346# bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[1] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3646 vdd dac_3v_8bit_0/b4a dac_3v_8bit_0/b4b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3647 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3648 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3649 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3650 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbp dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3651 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3652 dac_3v_column_odd_0[1].res_in0 dac_3v_column_odd_0[1].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3653 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3654 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output7.A a_n53197_n19329# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3655 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3656 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3657 a_30098_n21083# a_31605_n21083# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3658 dac_3v_column_odd_0[2].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_odd_0[2].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3659 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3660 dac_3v_column_odd_0[4].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_odd_0[4].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3661 dac_3v_column_0[2].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[2].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3662 a_25384_n14015# dac_3v_8bit_0/b0b dac_3v_column_0[5].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3663 dac_3v_column_odd_0[3].res_in0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[3].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=500000u
X3664 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n53615_n20961# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3665 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbp2 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3666 a_23170_n12950# dac_3v_8bit_0/b1a dac_3v_column_odd_0[4].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3667 a_22370_n8686# dac_3v_8bit_0/b0a dac_3v_column_odd_0[2].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3668 dac_3v_column_odd_0[2].res_in1 a_22370_n8686# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3669 a_n55858_5903# dvdd dvss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X3670 dvss dac_3v_8bit_0/b3a dac_3v_8bit_0/b3b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3671 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3672 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3673 dac_3v_8bit_0/b5a level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3674 a_26891_n9751# dac_3v_8bit_0/b0a dac_3v_column_0[3].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3675 a_n55794_10065# a_n55794_10065# a_n55858_8035# dvdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=1e+06u
X3676 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3677 dac_3v_8bit_0/b3a level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3678 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3679 a_22563_n13623# a_24070_n13623# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3680 dvdd bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3681 dac_3v_column_odd_0[6].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_odd_0[6].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3682 dvss a_27058_3107# a_27998_3404# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X3683 vdd level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3684 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3685 dac_3v_column_odd_0[0].dum_out1 vss a_34426_n5921# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3686 dac_3v_column_0[6].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_0[6].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3687 dac_3v_column_0[3].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_0[3].res1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3688 dvss bias_0.bi__pmirr_0.gate_cas dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3689 dac_3v_column_odd_0[6].out1_0_3 dac_3v_8bit_0/b0b a_31605_n17887# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3690 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3691 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.X a_n54945_n17689# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3692 dvss a_n55353_n19355# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3693 dac_3v_column_0[7].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_0[7].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3694 a_20863_n16581# vss a_20863_n16581# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3695 dac_3v_column_0[4].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[4].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3696 a_33719_n4698# vss dac_3v_column_odd_0[0].res_out1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3697 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3698 dac_3v_column_odd_0[2].out1_0_2 dac_3v_8bit_0/b0a a_28591_n9359# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3699 dac_3v_column_0[5].out0_2 dac_3v_8bit_0/b3a dac_3v_column_0[5].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X3700 dac_3v_column_odd_0[3].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[3].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3701 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3702 a_26891_n12950# a_28398_n12950# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3703 dvss level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b3a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3704 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3705 dvss dac_3v_8bit_0/b7b dac_3v_8bit_0/b7a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3706 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X3707 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3708 a_31412_n20410# vss a_31412_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3709 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3710 a_28591_n4028# a_30098_n4028# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3711 a_25384_n5487# dac_3v_8bit_0/b0b dac_3v_column_0[1].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3712 a_27084_n9359# a_28591_n9359# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3713 a_34426_n8053# vdd a_34426_n8053# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3714 dac_3v_column_odd_0[1].res_in1 vss a_20863_n6988# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X3715 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3716 vdd level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b1a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3717 a_31412_n15082# dac_3v_8bit_0/b0a dac_3v_column_odd_0[5].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3718 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3719 dac_3v_column_0[7].out1_0_2 dac_3v_8bit_0/b0a a_27084_n18952# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3720 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3721 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3722 a_31942_2371# a_31942_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3723 a_32919_n2724# vss a_32919_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3724 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3725 dac_3v_column_0[3].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[3].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3726 dac_3v_column_0[0].out1_0_3 dac_3v_8bit_0/b0a a_30098_n4028# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3727 dac_3v_column_odd_0[4].res_in0 dac_3v_column_odd_0[4].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3728 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3729 a_23170_n8686# dac_3v_8bit_0/b1b dac_3v_column_odd_0[2].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3730 a_23170_n4422# dac_3v_8bit_0/b1a dac_3v_column_odd_0[0].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3731 dac_3v_column_0[4].out1_0_1 dac_3v_8bit_0/b0b a_24070_n12556# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3732 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3733 dac_3v_column_odd_0[2].out1_0_3 dac_3v_8bit_0/b0a a_31605_n9359# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3734 dac_3v_column_0[2].res1_in a_22563_n8292# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3735 a_27691_n20686# vss a_27691_n20686# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3736 dac_3v_column_0[4].res1_in a_22370_n11883# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3737 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbn dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3738 dac_3v_column_0[0].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_0[0].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3739 a_31412_n14015# dac_3v_column_odd_0[4].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3740 dac_3v_column_0[2].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_0[2].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3741 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3742 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3743 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3744 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3745 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X3746 a_n55527_n18241# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n55599_n18241# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3747 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3748 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3749 dac_3v_column_odd_0[6].out4 dac_3v_8bit_0/b4b dac_3v_column_0[6].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3750 dvss level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b4a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3751 a_23877_n2724# vss a_23877_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3752 dac_3v_column_odd_0[4].out1_2 dac_3v_8bit_0/b2a dac_3v_column_odd_0[4].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3753 a_n54427_5925# bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__res_xhigh_po w=350000u l=7e+06u
X3754 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3755 a_31605_n4028# dac_3v_column_odd_0[0].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3756 dac_3v_column_0[5].res1_in vdd a_20863_n14449# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X3757 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3758 level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3759 a_29905_n5487# dac_3v_8bit_0/b0a dac_3v_column_0[1].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3760 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3761 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B a_n55353_n19355# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3762 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3763 dvss dac_3v_8bit_0/b6b dac_3v_8bit_0/b6a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3764 dac_3v_column_0[1].out1_0_2 dac_3v_8bit_0/b0a a_28591_n6160# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3765 a_20156_n6830# vdd a_20156_n6830# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+11p pd=7.74e+06u as=0p ps=0u w=1e+06u l=500000u
X3766 dac_3v_column_odd_0[0].out1_0_2 dac_3v_8bit_0/b0b a_28591_n5095# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3767 dac_3v_column_odd_0[2].out1_0_0 dac_3v_8bit_0/b0a a_22563_n9359# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3768 level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3769 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3770 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3771 dac_3v_column_0[6].out1_0_2 dac_3v_8bit_0/b0b a_28591_n16820# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3772 dac_3v_column_0[5].out_3 dac_3v_8bit_0/b3b dac_3v_column_0[5].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3773 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X3774 dac_3v_column_0[5].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_0[5].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3775 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3776 dac_3v_8bit_0/b5a level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3777 a_22563_n4028# a_24070_n4028# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3778 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3779 dac_3v_column_odd_0[5].out1_0_3 dac_3v_8bit_0/b0a a_31605_n15755# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3780 dac_3v_column_odd_0[4].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[4].res_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X3781 a_31412_n11883# dac_3v_8bit_0/b0a dac_3v_column_0[4].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3782 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3783 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3784 a_20156_n11094# vss a_20156_n11094# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3785 a_n48347_n15278# a_n48623_n15278# dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X3786 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3787 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3788 a_n25087_n925# a_n24701_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X3789 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3790 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3791 dvdd a_n54945_n17689# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.X dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3792 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3793 a_n54945_n21255# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3794 dac_3v_column_odd_0[0].out_5 dac_3v_8bit_0/b5b dac_3v_column_odd_0[0].out4 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3795 dac_3v_column_0[0].out1_0_1 dac_3v_8bit_0/b0b a_25577_n4028# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3796 dac_3v_column_0[1].out1_0_3 dac_3v_8bit_0/b0a a_31605_n6160# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3797 dvss dvss bandgap_0.bg__pnp_group_0.eg sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=1
X3798 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3799 a_24070_n18952# a_25577_n18952# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3800 a_n21740_n3691# bias_0.bi__amplifier_0.inn dvss dvss sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X3801 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._17_.X a_n55405_n20961# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3802 dvdd testbuffer_0.tb__mux_0.tbm__passgate_5.en a_n48623_n21248# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X3803 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X3804 dac_3v_column_odd_0[4].res_out1 dac_3v_8bit_0/b0b dac_3v_column_0[5].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X3805 a_25577_n20019# a_27084_n20019# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3806 vdd dac_3v_8bit_0/b6b dac_3v_8bit_0/b6a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3807 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3808 dvss level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3809 dac_3v_8bit_0/b2a level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3810 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3811 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X3812 dac_3v_column_0[1].out1_0_0 dac_3v_8bit_0/b0a a_22563_n6160# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3813 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3814 dac_3v_column_odd_0[6].out1_0_2 dac_3v_8bit_0/b0a a_28591_n17887# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3815 a_29905_n2290# vdd a_29905_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3816 dac_3v_column_0[7].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[7].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3817 a_25384_n17214# a_26891_n17214# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3818 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3819 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3820 dac_3v_8bit_0/b6a dac_3v_8bit_0/b6b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3821 a_34426_n14449# vss a_34426_n14449# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3822 a_33719_n13226# vdd dac_3v_column_odd_0[4].res_out1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3823 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3824 dac_3v_column_0[5].out0_1_0 dac_3v_8bit_0/b2a dac_3v_column_0[5].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3825 dac_3v_column_0[5].out0_1_1 dac_3v_8bit_0/b2a dac_3v_column_0[5].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3826 bias_0.bi__amplifier_0.mirr bias_0.bi__amplifier_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X3827 a_27084_n17887# a_28591_n17887# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3828 dac_3v_column_0[2].out0_1_1 dac_3v_8bit_0/b2a dac_3v_column_0[2].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3829 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3830 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._07_.X a_n55313_n22049# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3831 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3832 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3833 level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3834 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3835 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X3836 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3837 a_31412_n12950# dac_3v_8bit_0/b0b dac_3v_column_odd_0[4].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3838 a_22174_2371# a_22174_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3839 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3840 a_20156_n16423# vss dac_3v_column_0[6].dum1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3841 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3842 a_25384_n4422# a_26891_n4422# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3843 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3844 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3845 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X3846 testbuffer_0.tb__mux_0.tbm__passgate_4.en a_n55233_n20443# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3847 dac_3v_column_odd_0[3].out1_0_0 dac_3v_8bit_0/b0a a_22563_n11491# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3848 a_20863_n6988# vss a_20863_n6988# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3849 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3850 dac_3v_column_odd_0[5].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_odd_0[5].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3851 a_29264_2837# a_29626_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3852 vdd dac_3v_8bit_0/b3a dac_3v_8bit_0/b3b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3853 dac_3v_column_odd_0[3].out_3 dac_3v_8bit_0/b3a dac_3v_column_odd_0[3].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3854 dac_3v_column_odd_0[6].res_out1 dac_3v_column_odd_0[6].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3855 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3856 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3857 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._11_.A a_n55547_n19873# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3858 a_32919_n2290# vdd a_34426_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3859 a_n55646_9265# a_n55646_9265# a_n55794_10065# dvdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+11p pd=1.58e+06u as=0p ps=0u w=500000u l=1e+06u
X3860 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3861 a_23170_n19346# dac_3v_8bit_0/b1b dac_3v_column_odd_0[7].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3862 dac_3v_column_odd_0[4].out0_2 dac_3v_8bit_0/b3b dac_3v_column_odd_0[4].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3863 a_26891_n19346# dac_3v_8bit_0/b0a dac_3v_column_odd_0[7].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3864 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3865 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3866 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3867 dac_3v_8bit_0/b7b level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3868 dac_3v_column_odd_0[4].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[4].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3869 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3870 dvss a_29626_3404# a_29264_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3871 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3872 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3873 dvss dac_3v_8bit_0/b0b dac_3v_8bit_0/b0a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3874 a_25384_n2290# vdd a_25384_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3875 dvss level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b6b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3876 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3877 a_20156_n7895# vss dac_3v_column_0[2].dum1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X3878 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3879 dac_3v_8bit_0/b3b dac_3v_8bit_0/b3a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3880 a_23802_2206# a_23802_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X3881 a_20156_n6830# vdd dac_3v_column_odd_0[1].dum_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3882 dac_3v_column_odd_0[6].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_odd_0[6].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3883 a_20156_n17490# vdd dac_3v_column_odd_0[6].dum_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3884 a_28398_n8686# a_29905_n8686# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3885 vdd level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3886 dac_3v_column_odd_0[6].out1_2 dac_3v_8bit_0/b2b dac_3v_column_odd_0[6].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3887 a_25384_n18279# dac_3v_8bit_0/b0a dac_3v_column_0[7].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3888 dac_3v_8bit_0/b7a dac_3v_8bit_0/b7b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3889 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bias_basis_current_0.bb__nmirr_0.ibn bias_basis_current_0.bb__nmirr_0.ibn dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3890 dac_3v_column_0[7].res1_in vss a_20863_n18713# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3891 dac_3v_column_odd_0[7].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[7].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3892 dac_3v_column_0[3].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_0[3].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3893 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3894 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3895 a_31412_n10818# dac_3v_column_odd_0[3].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3896 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3897 level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3898 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3899 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3900 a_23170_n17214# dac_3v_8bit_0/b2b dac_3v_column_odd_0[6].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3901 a_n32750_n605# a_n31275_n477# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X3902 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3903 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3904 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3905 a_28591_n16820# a_30098_n16820# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3906 sbamuxm4_0/ibp[2] bias_0.bi__pmirr_0.gate a_n42353_12343# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3907 a_n25473_n925# a_n25859_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X3908 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output6.A a_n55047_n18669# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3909 dvss in[1] a_n55547_n19873# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3910 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3911 dvdd a_n54301_n18241# testbuffer_0.tb__mux_0.tbm__passgate_3.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3912 dac_3v_column_0[4].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[4].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3913 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3914 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3915 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3916 dac_3v_column_0[5].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_0[5].res1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3917 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3918 dvdd bias_0.bi__pmirr_0.gate a_n40589_12119# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X3919 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3920 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3921 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output8.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3922 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3923 dvss a_34510_3404# a_34148_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3924 dac_3v_column_odd_0[2].res_in0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[2].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3925 a_31412_n8686# dac_3v_column_odd_0[2].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3926 a_28398_n6554# dac_3v_8bit_0/b0b dac_3v_column_odd_0[1].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3927 vhigh dac_3v_column_0[0].dum0_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3928 dac_3v_column_0[1].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_0[1].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3929 dvss a_n53983_n17697# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3930 testbuffer_0.tb__mux_0.tbm__decoder3to8_0._21_.A a_n55681_n18241# dvss dvss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3931 a_n54400_n21689# a_n54587_n22049# a_n54487_n21933# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X3932 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3933 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3934 a_27084_n2963# a_28591_n2963# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3935 dac_3v_column_0[3].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_0[3].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3936 a_33719_n8962# vdd a_33719_n8962# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3937 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3938 dvdd bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3939 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3940 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3941 dac_3v_column_0[1].res1_in a_22370_n5487# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3942 a_22370_n5487# dac_3v_8bit_0/b0a dac_3v_column_0[1].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3943 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3944 a_28591_n8292# a_30098_n8292# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3945 vdd dac_3v_8bit_0/b5a dac_3v_8bit_0/b5b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3946 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3947 a_33719_n13226# vss dac_3v_column_odd_0[4].res_out1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3948 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3949 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X3950 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3951 dac_3v_column_odd_0[6].res_out1 dac_3v_8bit_0/b0a dac_3v_column_0[7].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3952 a_23877_n8686# dac_3v_8bit_0/b0b dac_3v_column_odd_0[2].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3953 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X3954 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3955 a_22563_n10424# a_24070_n10424# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3956 a_22370_n8686# a_23877_n8686# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3957 a_23877_n19346# a_25384_n19346# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3958 dac_3v_column_0[5].out0_1_0 dac_3v_8bit_0/b2b dac_3v_column_0[5].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3959 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3960 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3961 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3962 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3963 dvss a_n53523_n22049# testbuffer_0.tb__mux_0.tbm__passgate_5.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3964 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3965 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3966 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3967 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3968 a_23170_n8686# dac_3v_8bit_0/b2b dac_3v_column_odd_0[2].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3969 a_31412_n6554# dac_3v_8bit_0/b0b dac_3v_column_odd_0[1].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3970 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3971 testbuffer_0.tb__mux_0.tbm__passgate_2.en a_n53197_n19329# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3972 a_22370_n20844# vdd a_22370_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3973 dac_3v_column_0[7].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[7].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3974 sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X3975 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3976 a_34426_n11252# vdd a_34426_n11252# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3977 vdd level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b2a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3978 a_27084_n6160# a_28591_n6160# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3979 sbamuxm4_0/ibn[0] bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[0] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X3980 dac_3v_column_0[0].res1_in vss a_20863_n3789# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3981 a_n21999_n925# a_n22385_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X3982 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3983 dvss a_31942_3107# a_31942_2371# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3984 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3985 a_31605_n8292# dac_3v_column_odd_0[2].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3986 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3987 a_n55047_n18669# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvss dvss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X3988 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output8.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3989 dac_3v_column_odd_0[0].out4 dac_3v_8bit_0/b4a dac_3v_column_0[0].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3990 a_22370_n6554# dac_3v_8bit_0/b0b dac_3v_column_odd_0[1].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X3991 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3992 dac_3v_column_odd_0[7].dum_in0 vdd a_34426_n19780# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X3993 a_23170_n15082# dac_3v_8bit_0/b1a dac_3v_column_odd_0[5].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3994 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3995 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3996 dac_3v_column_0[6].dum1_in dac_3v_column_0[6].res1_in vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X3997 a_34426_n2724# vss a_34426_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3998 dac_3v_column_0[1].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[1].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X3999 a_n46909_n24233# a_n47185_n24233# dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X4000 a_33719_n3631# vdd dac_3v_column_odd_0[0].res_in0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4001 dac_3v_column_odd_0[2].out0_2 dac_3v_8bit_0/b3b dac_3v_column_odd_0[2].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4002 dac_3v_8bit_0/b6a dac_3v_8bit_0/b6b vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4003 a_23170_n4422# dac_3v_8bit_0/b2a dac_3v_column_odd_0[0].out0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4004 dac_3v_column_odd_0[1].res_out1 dac_3v_8bit_0/b0a dac_3v_column_0[2].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=500000u
X4005 dvss dvss bandgap_0.bg__pnp_group_0.eg sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=1
X4006 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4007 dac_3v_column_odd_0[3].out1_0_1 dac_3v_8bit_0/b0b a_25577_n11491# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X4008 a_22563_n8292# a_24070_n8292# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4009 dac_3v_8bit_0/b6b level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4010 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4011 dvss a_n53197_n22593# testbuffer_0.tb__mux_0.tbm__passgate_7.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4012 dac_3v_column_0[2].out_3 dac_3v_8bit_0/b3b dac_3v_column_0[2].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4013 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4014 dvss dac_3v_8bit_0/b2a dac_3v_8bit_0/b2b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4015 dac_3v_column_0[0].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[0].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4016 a_23877_n16147# a_25384_n16147# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4017 level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4018 dvss level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4019 dac_3v_column_0[3].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[3].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4020 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._16_.C a_n54440_n20729# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.0785e+11p ps=1.36e+06u w=420000u l=150000u
X4021 vdd dac_3v_8bit_0/b6b dac_3v_8bit_0/b6a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4022 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X4023 a_25384_n2724# vss a_25384_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4024 a_23170_n19346# dac_3v_8bit_0/b1b dac_3v_column_odd_0[7].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4025 testbuffer_0.tb__mux_0.tbm__passgate_5.en a_n53523_n22049# dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4026 a_n32750_2575# a_n31275_2703# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X4027 a_20156_n3631# vdd a_20156_n3631# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4028 dac_3v_column_0[2].out1_0_2 dac_3v_8bit_0/b0b a_27084_n8292# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4029 dac_3v_column_0[0].out1_0_1 dac_3v_8bit_0/b0b a_24070_n4028# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4030 a_26008_2837# a_26370_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4031 a_20156_n2566# vss a_20156_n2566# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4032 a_23877_n7619# dac_3v_8bit_0/b0a dac_3v_column_0[2].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4033 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4034 dvss dac_3v_8bit_0/b5a dac_3v_8bit_0/b5b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4035 dac_3v_column_odd_0[0].out1_0_3 dac_3v_8bit_0/b0b a_30098_n5095# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4036 a_28398_n20410# a_29905_n20410# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4037 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4038 a_20863_n4856# vdd a_20863_n4856# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4039 dac_3v_column_0[4].out1_0_3 dac_3v_8bit_0/b0a a_31605_n12556# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4040 dac_3v_column_0[3].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_0[3].res1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4041 sbamuxm4_0/vb[0] a_n32029_12624# dvss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X4042 dvss bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4043 dvss a_26370_3404# a_26008_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4044 dac_3v_8bit_0/b3b dac_3v_8bit_0/b3a vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4045 a_11923_n7894# a_17355_n7576# vss sky130_fd_pr__res_xhigh_po w=350000u l=2.5e+07u
X4046 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4047 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X4048 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4049 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4050 dac_3v_column_odd_0[6].out1_0_0 dac_3v_8bit_0/b0b a_22563_n17887# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X4051 dac_3v_column_0[7].out1_0_1 dac_3v_8bit_0/b1a dac_3v_column_0[7].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4052 dac_3v_column_0[4].out0_1_1 dac_3v_8bit_0/b1a dac_3v_column_0[4].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4053 dvss level_shifter_array_0/level_shifter_0[4].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b4a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4054 dvdd bias_0.bi__pmirr_0.gate dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X4055 dvss dac_3v_8bit_0/b2a dac_3v_8bit_0/b2b dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4056 a_20156_n18555# vss a_20156_n18555# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4057 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4058 dac_3v_column_odd_0[0].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_odd_0[0].res_in1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4059 a_29905_n2724# vss a_29905_n2724# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4060 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4061 vdd level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b7b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4062 dac_3v_column_0[0].out1_0_2 dac_3v_8bit_0/b0a a_27084_n4028# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X4063 a_25384_n20410# vss a_25384_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4064 dac_3v_column_odd_0[1].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_odd_0[1].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4065 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4066 dvdd a_n53197_n22593# testbuffer_0.tb__mux_0.tbm__passgate_7.en dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4067 a_25384_n15082# dac_3v_8bit_0/b0a dac_3v_column_odd_0[5].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X4068 dac_3v_column_0[7].out1_0_2 dac_3v_8bit_0/b0b a_27084_n18952# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4069 dac_3v_column_odd_0[5].res_in1 vss a_20863_n15516# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.655e+11p ps=5.64e+06u w=650000u l=500000u
X4070 dvss testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output4.A dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4071 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4072 a_n32750_n2725# a_n31275_n2597# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X4073 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4074 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A a_n53645_n19873# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4075 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4076 dac_3v_8bit_0/b3a level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4077 dvdd testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4078 dac_3v_column_odd_0[2].dum_in1 dac_3v_column_odd_0[2].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4079 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X4080 a_27691_n20686# vdd a_27691_n20686# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4081 dvdd a_n53983_n17697# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._10_.X dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4082 dac_3v_column_odd_0[7].out_3 dac_3v_8bit_0/b3b dac_3v_column_odd_0[7].out1_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4083 a_28591_n13623# a_30098_n13623# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4084 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbn2 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4085 dac_3v_column_odd_0[7].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[7].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4086 a_25384_n14015# a_26891_n14015# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4087 a_33719_n10027# vdd dac_3v_column_odd_0[3].res_in0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4088 bandgap_0.bg__pnp_group_0.eg dvss a_n31275_583# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X4089 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4090 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4091 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4092 vdd level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4093 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4094 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4095 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_0.diffb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4096 a_27058_2371# a_27058_3107# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4097 a_27084_n14688# a_28591_n14688# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4098 dac_3v_column_odd_0[1].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_odd_0[1].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4099 a_22370_n10818# dac_3v_8bit_0/b0a dac_3v_column_odd_0[3].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X4100 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd10 bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.mirr dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X4101 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4102 a_29905_n17214# dac_3v_8bit_0/b0a dac_3v_column_odd_0[6].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4103 bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__pmirr_0.vbp dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4104 sbamuxm4_0/ibn[1] bias_0.bi__pmirr_0.gate_cas sbamuxm4_0/ibn[1] dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4105 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4106 bias_0.bi__amplifier_0.mirr bias_0.bi__amplifier_0.mirr dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X4107 vdd level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b0b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4108 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4109 a_31605_n18952# dac_3v_column_odd_0[7].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4110 a_20024_n21083# a_20863_n20410# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4111 level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_4_0.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4112 testbuffer_0.tb__mux_0.tbm__passgate_2.out a_n47185_n18263# inp[3] dvdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4113 dvss a_29626_3404# a_29264_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4114 a_n53983_n17697# testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4115 vdd dac_3v_8bit_0/b1a dac_3v_8bit_0/b1b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4116 a_20863_n2290# a_22370_n2290# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4117 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4118 bias_basis_current_0.bb__pmirr_0.vbp bias_basis_current_0.bb__pmirr_0.vbn bias_basis_current_0.bb__nmirr_0.vres dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4119 a_34148_2837# a_34510_3404# dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4120 a_20863_n18713# vdd a_20863_n18713# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4121 a_20863_n20410# a_22563_n21083# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4122 dac_3v_column_0[4].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_0[4].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4123 dac_3v_column_odd_0[5].res_in0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[5].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4124 dac_3v_column_odd_0[1].out1_0_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[1].out1_1_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4125 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4126 dac_3v_8bit_0/b3a level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4127 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4128 dac_3v_column_odd_0[5].res_in0 dac_3v_column_odd_0[5].dum_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4129 a_25384_n11883# dac_3v_8bit_0/b0a dac_3v_column_0[4].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X4130 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4131 dvdd a_33570_3107# a_34510_3404# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X4132 dac_3v_8bit_0/b7a dac_3v_8bit_0/b7b dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4133 dac_3v_column_odd_0[5].out1_0_1 dac_3v_8bit_0/b0a a_25577_n15755# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4134 a_29905_n9751# dac_3v_8bit_0/b0b dac_3v_column_0[3].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X4135 dac_3v_column_0[4].res1_in vss a_20863_n12317# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4136 dac_3v_column_0[6].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[6].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4137 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4138 a_22370_n15082# a_23877_n15082# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4139 dac_3v_column_odd_0[3].out1_0_3 dac_3v_8bit_0/b0b a_31605_n11491# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X4140 a_26891_n16147# dac_3v_8bit_0/b0a dac_3v_column_0[6].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4141 dvss bias_0.bi__pmirr_0.gate_cas dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4142 dvss a_30314_3107# a_31254_3404# dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X4143 a_20863_n20410# vdd a_20863_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4144 dac_3v_column_0[3].out1_2 dac_3v_8bit_0/b2b dac_3v_column_0[3].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4145 dvss a_n54301_n18241# testbuffer_0.tb__mux_0.tbm__passgate_3.en dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4146 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4147 a_34426_n19780# vss a_34426_n19780# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4148 dvdd bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X4149 dac_3v_column_odd_0[7].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[7].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4150 dac_3v_column_odd_0[5].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[5].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4151 a_33719_n6830# vss a_33719_n6830# vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.655e+11p pd=5.64e+06u as=0p ps=0u w=650000u l=500000u
X4152 a_26891_n2290# vdd a_26891_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X4153 a_26891_n20844# vdd a_26891_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4154 a_n23157_n925# a_n22771_2107# dvss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X4155 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X4156 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4157 a_22370_n20844# vss a_22370_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4158 dac_3v_column_0[2].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_0[2].res1_in vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4159 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4160 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4161 a_28398_n5487# a_29905_n5487# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4162 a_23877_n6554# a_25384_n6554# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4163 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4164 dvdd a_n55353_n19355# testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.B dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4165 dac_3v_column_odd_0[2].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_odd_0[2].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4166 dac_3v_column_odd_0[1].res_out1 dac_3v_column_odd_0[1].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4167 a_25430_2206# a_25430_2371# vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X4168 a_27691_n2566# vdd a_27691_n2566# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4169 a_30098_n15755# a_31605_n15755# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4170 dac_3v_column_odd_0[4].dum_in1 dac_3v_column_odd_0[4].res_in1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4171 dac_3v_column_odd_0[2].dum_out1 vdd a_34426_n10185# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X4172 testbuffer_0.tb__mux_0.tbm__decoder3to8_0.output6.A testbuffer_0.tb__mux_0.tbm__decoder3to8_0._20_.A dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4173 dac_3v_column_0[6].out1_0_0 dac_3v_8bit_0/b1a dac_3v_column_0[6].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4174 level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__inv_4_0.A level_shifter_array_0/level_shifter_0[7].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4175 dac_3v_column_odd_0[7].out4 dac_3v_8bit_0/b4a dac_3v_column_0[7].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4176 dac_3v_column_odd_0[0].res_in0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[0].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4177 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4178 dac_3v_column_0[5].out1_0_2 dac_3v_8bit_0/b1b dac_3v_column_0[5].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4179 dac_3v_8bit_0/b2a level_shifter_array_0/level_shifter_0[2].sky130_fd_sc_hvl__inv_8_1.A vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4180 dac_3v_column_odd_0[3].res_out1 dac_3v_8bit_0/b0a dac_3v_column_0[4].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4181 dac_3v_column_0[5].out0_1_1 dac_3v_8bit_0/b2b dac_3v_column_0[5].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4182 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4183 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4184 vdd level_shifter_array_0/level_shifter_0[3].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b3a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4185 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4186 a_23877_n12950# a_25384_n12950# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4187 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4188 dvss bias_0.bi__amplifier_0.bias bias_0.bi__amplifier_0.bias dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X4189 bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.diff bandgap_0.bg__se_folded_cascode_p_0.bgfc__pmirr_0.vbp1 dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4190 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4191 vlow vdd a_32919_n20844# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4192 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4193 a_25384_n9751# dac_3v_8bit_0/b0a dac_3v_column_0[3].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X4194 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4195 dvss a_23114_3404# a_22752_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4196 a_25384_n12950# dac_3v_8bit_0/b0b dac_3v_column_odd_0[4].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4197 dvdd bias_0.bi__pmirr_0.gate a_n40589_11895# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X4198 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X4199 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4200 a_26891_n8686# dac_3v_8bit_0/b0a dac_3v_column_odd_0[2].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4201 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4202 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.mirr sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X4203 a_28398_n3355# dac_3v_8bit_0/b0b dac_3v_column_0[0].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4204 a_23877_n4422# dac_3v_8bit_0/b0a dac_3v_column_odd_0[0].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4205 a_31412_n5487# dac_3v_column_odd_0[0].res_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4206 dac_3v_column_odd_0[0].res_out1 dac_3v_8bit_0/b0b dac_3v_column_0[1].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4207 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4208 dac_3v_8bit_0/b5b dac_3v_8bit_0/b5a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4209 dac_3v_column_0[7].out1_0_3 dac_3v_8bit_0/b0b a_30098_n18952# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4210 dac_3v_column_odd_0[2].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_odd_0[2].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4211 dvss testbuffer_0.tb__mux_0.tbm__passgate_1.en a_n48623_n15278# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X4212 dac_3v_column_0[7].out1_0_1 dac_3v_8bit_0/b0a a_24070_n18952# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X4213 vdd follower_amp_0.pdrv2 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4214 vdd level_shifter_array_0/level_shifter_0[6].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b6b vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4215 dac_3v_column_odd_0[5].out1_0_1 dac_3v_8bit_0/b1b dac_3v_column_odd_0[5].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4216 dac_3v_column_0[4].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_0[4].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4217 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X4218 dac_3v_8bit_0/b2b dac_3v_8bit_0/b2a dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4219 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4220 a_34426_n20844# vss a_34426_n20844# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4221 a_20863_n15516# vss a_20863_n15516# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4222 a_33719_n5763# vdd a_33719_n5763# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4223 dac_3v_column_odd_0[6].out1_0_3 dac_3v_8bit_0/b1a dac_3v_column_odd_0[6].out1_1_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4224 vdd level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4225 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4226 dac_3v_column_odd_0[1].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[1].out0_0_1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4227 dvss dvss bandgap_0.bg__pnp_group_0.eg sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=1
X4228 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4229 a_30705_n20686# vdd a_30705_n20686# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4230 dac_3v_column_odd_0[4].out0_2 dac_3v_8bit_0/b3a dac_3v_column_odd_0[4].out_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4231 bias_0.bi__pmirr_0.gate bias_0.bi__pmirr_0.fb sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X4232 a_24677_n20686# vss a_24677_n20686# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4233 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X4234 a_33719_n10027# vss dac_3v_column_odd_0[3].res_in0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4235 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p sbamuxm4_0/ibp[0] testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__cascode_p_0.outs1 dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X4236 a_23877_n5487# dac_3v_8bit_0/b0b dac_3v_column_0[1].out0_0_3 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X4237 dac_3v_column_0[1].out1_0_2 dac_3v_8bit_0/b1a dac_3v_column_0[1].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4238 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1n bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4239 dvss dvss dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4240 a_22370_n5487# a_23877_n5487# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4241 dvss level_shifter_array_0/level_shifter_0[1].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b1a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4242 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4243 dac_3v_column_odd_0[6].out0_1_0 dac_3v_8bit_0/b1a dac_3v_column_odd_0[6].out0_0_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4244 a_20156_n15358# vss a_20156_n15358# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4245 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4246 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X4247 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4248 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out dvss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4249 dvss level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__inv_8_1.A dac_3v_8bit_0/b5a dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4250 dac_3v_column_odd_0[0].res_out1 dac_3v_column_odd_0[0].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4251 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4252 a_31412_n3355# dac_3v_8bit_0/b0b dac_3v_column_0[0].out0_0_0 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4253 dac_3v_column_0[1].out0_1_1 dac_3v_8bit_0/b2b dac_3v_column_0[1].out0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4254 bias_0.bi__amplifier_0.bias bias_0.bi__amplifier_0.bias dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X4255 vss follower_amp_0.ndrv dac_out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4256 dac_3v_column_odd_0[6].out1_0_2 dac_3v_8bit_0/b0a a_27084_n17887# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X4257 a_23170_n8686# dac_3v_8bit_0/b1a dac_3v_column_odd_0[2].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4258 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4259 a_30705_n2566# vss a_30098_n2963# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X4260 dac_3v_column_odd_0[7].out1_0_0 dac_3v_8bit_0/b0a dac_3v_column_odd_0[7].res_in1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4261 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1p testbuffer_0.tb__mux_0.tbm__passgate_2.out testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4262 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4263 a_23802_3107# b6 dvss dvss sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X4264 dac_3v_column_0[5].out1_2 dac_3v_8bit_0/b2a dac_3v_column_0[5].out1_1_0 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4265 a_22370_n2724# vdd a_22370_n2724# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4266 dac_3v_column_odd_0[3].out1_0_2 dac_3v_8bit_0/b0a a_28591_n11491# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4267 vdd dac_3v_8bit_0/b0b dac_3v_8bit_0/b0a vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4268 a_22370_n3355# dac_3v_8bit_0/b0b dac_3v_column_0[0].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4269 dac_out follower_amp_0.ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4270 a_n46909_n15278# a_n47185_n15278# dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X4271 dvss testbuffer_0.tb__mux_0.tbm__passgate_2.en a_n47185_n18263# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X4272 dac_3v_column_0[0].out_3 dac_3v_8bit_0/b3a dac_3v_column_0[0].out1_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4273 dac_3v_column_0[1].out1_0_3 dac_3v_8bit_0/b1b dac_3v_column_0[1].out1_1_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4274 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X4275 dvss dvdd dvss dvss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X4276 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1p dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4277 dac_out follower_amp_0.pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4278 dac_3v_column_odd_0[5].dum_out1 vdd a_34426_n16581# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X4279 dac_3v_column_odd_0[5].out4 dac_3v_8bit_0/b4a dac_3v_column_odd_0[5].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4280 a_25384_n10818# a_26891_n10818# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4281 dvss testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.vbn1 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.outb1n dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4282 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4283 dac_3v_column_odd_0[7].out0_1_0 dac_3v_8bit_0/b1b dac_3v_column_odd_0[7].out0_0_1 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4284 dac_3v_column_odd_0[4].res_in1 vdd a_20863_n13384# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4285 sbamuxm4_0/ibn[0] bias_0.bi__pmirr_0.gate_cas a_n41084_7938# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4286 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out1p bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.vbn1 dvss dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4287 dvdd testbuffer_0.tb__mux_0.tbm__decoder3to8_0.input1.X a_n55681_n18241# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4288 a_31412_n19346# dac_3v_column_odd_0[7].res_in0 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4289 dac_3v_column_odd_0[0].out1_0_2 dac_3v_8bit_0/b0a a_28591_n5095# vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4290 dac_3v_column_0[1].out0_2 dac_3v_8bit_0/b3b dac_3v_column_0[1].out_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4291 vdd follower_amp_0.pdrv1 dac_out vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4292 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4293 a_27084_n11491# a_28591_n11491# vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
X4294 dac_3v_column_0[5].out1_0_0 dac_3v_8bit_0/b0b dac_3v_column_0[5].res1_in vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4295 bandgap_0.bg__se_folded_cascode_p_0.bgfc__casn_top_0.out bias_basis_current_0.bb__nmirr_0.ibn bandgap_0.bg__se_folded_cascode_p_0.bgfc__casp_top_0.nd11 dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X4296 dac_3v_column_odd_0[1].dum_out1 vss a_34426_n8053# vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4297 dac_out follower_amp_0.pdrv2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X4298 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4299 dvdd dvss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X4300 sbamuxm4_0/ibp[1] bias_0.bi__pmirr_0.gate a_n42353_11447# dvdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X4301 dvss bias_0.bi__nmirr_0.gate_n a_n42000_8994# dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X4302 a_20156_n12159# vss a_20156_n12159# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4303 dac_3v_column_odd_0[5].out1_0_2 dac_3v_8bit_0/b0b a_28591_n15755# vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.885e+11p ps=1.88e+06u w=650000u l=500000u
X4304 a_33719_n6830# vss dac_3v_column_odd_0[1].res_out1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4305 testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__pmirr_upper_0.outa1n sbamuxm4_0/muxout testbuffer_0.tb__se_folded_cascode_np_ab_0.tbfc__nmirr_0.diffa dvss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4306 dvss a_26370_3404# a_26008_2837# dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X4307 level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_8_1.A level_shifter_array_0/level_shifter_0[0].sky130_fd_sc_hvl__inv_4_0.A dvss dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4308 dvss a_25430_2206# level_shifter_array_0/level_shifter_0[5].sky130_fd_sc_hvl__lsbuflv2hv_1_0.X dvss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X4309 dac_3v_column_0[6].out0_1_1 dac_3v_8bit_0/b1b dac_3v_column_0[6].out0_0_2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4310 a_26891_n10818# dac_3v_8bit_0/b0b dac_3v_column_odd_0[3].out0_0_2 vdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X4311 a_22370_n10818# dac_3v_8bit_0/b0b dac_3v_column_odd_0[3].out0_0_3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.885e+11p pd=1.88e+06u as=0p ps=0u w=650000u l=500000u
X4312 dac_3v_column_odd_0[3].res_out1 dac_3v_column_odd_0[3].dum_out1 vss sky130_fd_pr__res_high_po w=350000u l=3e+06u
.ends

