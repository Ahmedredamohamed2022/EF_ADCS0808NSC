VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_ADCS0808NSC
  CLASS BLOCK ;
  FOREIGN EF_ADCS0808NSC ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END EF_ADCS0808NSC
END LIBRARY

